module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [18:0] __in0,
  output logic [14:0] __out0);
  logic [47:0] gzdLLzicase66426;
  logic [44:0] callRes;
  logic [47:0] gzdLLzicase66426R1;
  logic [44:0] callResR1;
  logic [47:0] gzdLLzicase66426R2;
  logic [44:0] callResR2;
  logic [47:0] gzdLLzicase66426R3;
  logic [44:0] callResR3;
  logic [47:0] gzdLLzicase66426R4;
  logic [44:0] callResR4;
  logic [47:0] gzdLLzicase66426R5;
  logic [44:0] callResR5;
  logic [47:0] gzdLLzicase66426R6;
  logic [44:0] callResR6;
  logic [47:0] gzdLLzicase66426R7;
  logic [44:0] callResR7;
  logic [47:0] gzdLLzicase66426R8;
  logic [44:0] callResR8;
  logic [47:0] gzdLLzicase66426R9;
  logic [44:0] callResR9;
  logic [47:0] gzdLLzicase66426R10;
  logic [44:0] callResR10;
  logic [47:0] gzdLLzicase66426R11;
  logic [44:0] callResR11;
  logic [0:0] __continue;
  logic [3:0] __resumption_tag;
  logic [24:0] __st0;
  logic [3:0] __resumption_tag_next;
  logic [24:0] __st0_next;
  assign gzdLLzicase66426 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426 (gzdLLzicase66426[43:19], gzdLLzicase66426[18:0], callRes);
  assign gzdLLzicase66426R1 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R1 (gzdLLzicase66426R1[43:19], gzdLLzicase66426R1[18:0], callResR1);
  assign gzdLLzicase66426R2 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R2 (gzdLLzicase66426R2[43:19], gzdLLzicase66426R2[18:0], callResR2);
  assign gzdLLzicase66426R3 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R3 (gzdLLzicase66426R3[43:19], gzdLLzicase66426R3[18:0], callResR3);
  assign gzdLLzicase66426R4 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R4 (gzdLLzicase66426R4[43:19], gzdLLzicase66426R4[18:0], callResR4);
  assign gzdLLzicase66426R5 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R5 (gzdLLzicase66426R5[43:19], gzdLLzicase66426R5[18:0], callResR5);
  assign gzdLLzicase66426R6 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R6 (gzdLLzicase66426R6[43:19], gzdLLzicase66426R6[18:0], callResR6);
  assign gzdLLzicase66426R7 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R7 (gzdLLzicase66426R7[43:19], gzdLLzicase66426R7[18:0], callResR7);
  assign gzdLLzicase66426R8 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R8 (gzdLLzicase66426R8[43:19], gzdLLzicase66426R8[18:0], callResR8);
  assign gzdLLzicase66426R9 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R9 (gzdLLzicase66426R9[43:19], gzdLLzicase66426R9[18:0], callResR9);
  assign gzdLLzicase66426R10 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R10 (gzdLLzicase66426R10[43:19], gzdLLzicase66426R10[18:0], callResR10);
  assign gzdLLzicase66426R11 = {{__resumption_tag, __st0}, __in0};
  zdLLzicase66426  zdLLzicase66426R11 (gzdLLzicase66426R11[43:19], gzdLLzicase66426R11[18:0], callResR11);
  assign {__continue, __out0, __resumption_tag_next, __st0_next} = (gzdLLzicase66426R11[47:44] == 4'h0) ? callResR11 : ((gzdLLzicase66426R10[47:44] == 4'h1) ? callResR10 : ((gzdLLzicase66426R9[47:44] == 4'h2) ? callResR9 : ((gzdLLzicase66426R8[47:44] == 4'h3) ? callResR8 : ((gzdLLzicase66426R7[47:44] == 4'h4) ? callResR7 : ((gzdLLzicase66426R6[47:44] == 4'h5) ? callResR6 : ((gzdLLzicase66426R5[47:44] == 4'h6) ? callResR5 : ((gzdLLzicase66426R4[47:44] == 4'h7) ? callResR4 : ((gzdLLzicase66426R3[47:44] == 4'h8) ? callResR3 : ((gzdLLzicase66426R2[47:44] == 4'h9) ? callResR2 : ((gzdLLzicase66426R1[47:44] == 4'ha) ? callResR1 : callRes))))))))));
  initial {__resumption_tag, __st0} <= 29'h0c000000;
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      {__resumption_tag, __st0} <= 29'h0c000000;
    end else begin
      {__resumption_tag, __st0} <= {__resumption_tag_next, __st0_next};
    end
  end
endmodule

module zdLLzicase62993 (input logic [0:0] arg0,
  input logic [0:0] arg1,
  input logic [0:0] arg2,
  input logic [0:0] arg3,
  input logic [0:0] arg4,
  input logic [0:0] arg5,
  input logic [0:0] arg6,
  input logic [0:0] arg7,
  input logic [0:0] arg8,
  input logic [0:0] arg9,
  input logic [0:0] arg10,
  input logic [0:0] arg11,
  input logic [0:0] arg12,
  input logic [0:0] arg13,
  input logic [0:0] arg14,
  input logic [0:0] arg15,
  input logic [0:0] arg16,
  input logic [0:0] arg17,
  input logic [0:0] arg18,
  input logic [0:0] arg19,
  input logic [0:0] arg20,
  input logic [0:0] arg21,
  input logic [2:0] arg22,
  output logic [24:0] res);
  assign res = {arg0, arg1, arg2, 1'h1, arg4, arg5, arg6, arg7, arg8, arg9, arg10, arg11, arg12, arg13, arg14, arg15, arg16, arg17, arg18, arg19, arg20, arg21, 3'h0};
endmodule

module zdLLzicase63071 (input logic [0:0] arg0,
  input logic [0:0] arg1,
  input logic [0:0] arg2,
  input logic [0:0] arg3,
  input logic [0:0] arg4,
  input logic [0:0] arg5,
  input logic [0:0] arg6,
  input logic [0:0] arg7,
  input logic [0:0] arg8,
  input logic [0:0] arg9,
  input logic [0:0] arg10,
  input logic [0:0] arg11,
  input logic [0:0] arg12,
  input logic [0:0] arg13,
  input logic [0:0] arg14,
  input logic [0:0] arg15,
  input logic [0:0] arg16,
  input logic [0:0] arg17,
  input logic [0:0] arg18,
  input logic [0:0] arg19,
  input logic [0:0] arg20,
  input logic [0:0] arg21,
  input logic [2:0] arg22,
  output logic [24:0] res);
  assign res = {arg0, arg1, arg2, 1'h1, arg4, arg5, arg6, arg7, arg8, arg9, arg10, arg11, arg12, arg13, arg14, 1'h1, arg16, arg17, arg18, arg19, arg20, arg21, 3'h0};
endmodule

module zdLLzicase63123 (input logic [0:0] arg0,
  input logic [0:0] arg1,
  input logic [0:0] arg2,
  input logic [0:0] arg3,
  input logic [0:0] arg4,
  input logic [0:0] arg5,
  input logic [0:0] arg6,
  input logic [0:0] arg7,
  input logic [0:0] arg8,
  input logic [0:0] arg9,
  input logic [0:0] arg10,
  input logic [0:0] arg11,
  input logic [0:0] arg12,
  input logic [0:0] arg13,
  input logic [0:0] arg14,
  input logic [0:0] arg15,
  input logic [0:0] arg16,
  input logic [0:0] arg17,
  input logic [0:0] arg18,
  input logic [0:0] arg19,
  input logic [0:0] arg20,
  input logic [0:0] arg21,
  input logic [2:0] arg22,
  output logic [24:0] res);
  assign res = {arg0, arg1, arg2, arg3, arg4, arg5, arg6, arg7, arg8, arg9, arg10, arg11, arg12, arg13, arg14, arg15, arg16, arg17, arg18, arg19, arg20, arg21, 3'h0};
endmodule

module zdLLzicase63392 (input logic [0:0] arg0,
  input logic [0:0] arg1,
  input logic [0:0] arg2,
  input logic [0:0] arg3,
  input logic [0:0] arg4,
  input logic [0:0] arg5,
  input logic [0:0] arg6,
  input logic [0:0] arg7,
  input logic [0:0] arg8,
  input logic [0:0] arg9,
  input logic [0:0] arg10,
  input logic [0:0] arg11,
  input logic [0:0] arg12,
  input logic [0:0] arg13,
  input logic [0:0] arg14,
  input logic [0:0] arg15,
  input logic [0:0] arg16,
  input logic [0:0] arg17,
  input logic [0:0] arg18,
  input logic [0:0] arg19,
  input logic [0:0] arg20,
  input logic [0:0] arg21,
  input logic [2:0] arg22,
  output logic [24:0] res);
  assign res = {arg0, arg1, 1'h1, arg3, arg4, arg5, arg6, arg7, arg8, arg9, arg10, arg11, arg12, arg13, arg14, arg15, arg16, arg17, arg18, arg19, arg20, arg21, arg22};
endmodule

module zdLLzicase63625 (input logic [0:0] arg0,
  input logic [0:0] arg1,
  input logic [0:0] arg2,
  input logic [0:0] arg3,
  input logic [0:0] arg4,
  input logic [0:0] arg5,
  input logic [0:0] arg6,
  input logic [0:0] arg7,
  input logic [0:0] arg8,
  input logic [0:0] arg9,
  input logic [0:0] arg10,
  input logic [0:0] arg11,
  input logic [0:0] arg12,
  input logic [0:0] arg13,
  input logic [0:0] arg14,
  input logic [0:0] arg15,
  input logic [0:0] arg16,
  input logic [0:0] arg17,
  input logic [0:0] arg18,
  input logic [0:0] arg19,
  input logic [0:0] arg20,
  input logic [0:0] arg21,
  input logic [2:0] arg22,
  output logic [24:0] res);
  assign res = {arg0, arg1, arg2, arg3, 1'h1, arg5, arg6, arg7, arg8, arg9, arg10, arg11, arg12, arg13, arg14, arg15, arg16, arg17, arg18, arg19, arg20, arg21, 3'h3};
endmodule

module zdLLzicase66426 (input logic [24:0] arg0,
  input logic [18:0] arg1,
  output logic [44:0] res);
  logic [43:0] gMainzidispatch;
  logic [49:0] gzdLLzilambda67585;
  logic [49:0] gzdLLzilambda62519;
  logic [24:0] gMainzilinkzustate;
  logic [24:0] gzdLLzicase62798;
  logic [27:0] gzdLLzilambda67580;
  logic [27:0] gzdLLzicase67578;
  logic [63:0] gzdLLzilambda67575;
  logic [63:0] gzdLLzicase67572;
  logic [46:0] gzdLLzilambda62558;
  logic [46:0] gzdLLzicase67541;
  logic [43:0] gzdLLzicase62545;
  logic [43:0] gMainzislsmzurun;
  logic [68:0] gzdLLzilambda67401;
  logic [68:0] gzdLLzicase67398;
  logic [68:0] gzdLLzilambda63819;
  logic [24:0] gzdLLzicase63730;
  logic [43:0] gzdLLzilambda67090;
  logic [43:0] gzdLLzicase67087;
  logic [43:0] gzdLLzilambda63816;
  logic [68:0] gzdLLzilambda67083;
  logic [68:0] gzdLLzicase67080;
  logic [68:0] gzdLLzilambda63813;
  logic [24:0] gMainzisendzutimezucode;
  logic [0:0] callRes;
  logic [44:0] gzdLLzilambda67076;
  logic [44:0] gzdLLzicase67073;
  logic [44:0] gzdLLzilambda63810;
  logic [69:0] gzdLLzilambda67069;
  logic [69:0] gzdLLzicase67065;
  logic [69:0] gzdLLzilambda63807;
  logic [25:0] gzdLLzicase63755;
  logic [0:0] gReWireziPreludezinot;
  logic [0:0] lit;
  logic [0:0] litR1;
  logic [43:0] gzdLLzilambda67060;
  logic [43:0] gzdLLzicase67057;
  logic [43:0] gzdLLzilambda63803;
  logic [68:0] gzdLLzilambda67053;
  logic [68:0] gzdLLzicase67050;
  logic [68:0] gzdLLzilambda63800;
  logic [24:0] gMainzilinkzudisablezuzz1;
  logic [0:0] callResR1;
  logic [44:0] gzdLLzilambda67046;
  logic [44:0] gzdLLzicase67043;
  logic [44:0] gzdLLzilambda63797;
  logic [69:0] gzdLLzilambda67039;
  logic [69:0] gzdLLzicase67035;
  logic [69:0] gzdLLzilambda63794;
  logic [24:0] gMainzirxzuerrorzusync;
  logic [0:0] callResR2;
  logic [45:0] gzdLLzilambda67030;
  logic [45:0] gzdLLzicase67026;
  logic [45:0] gzdLLzilambda63790;
  logic [1:0] gReWireziPreludezizbzb;
  logic [0:0] callResR3;
  logic [1:0] gReWireziPreludezizbzbR1;
  logic [0:0] callResR4;
  logic [25:0] id;
  logic [25:0] gzdLLzicase67021;
  logic [24:0] gzdLLzicase63783;
  logic [49:0] gzdLLzilambda66605;
  logic [49:0] gzdLLzilambda63781;
  logic [24:0] gzdLLzicase62993;
  logic [24:0] callResR5;
  logic [43:0] gzdLLzilambda67017;
  logic [43:0] gzdLLzicase66831;
  logic [39:0] callResR6;
  logic [39:0] gzdLLzilambda67428;
  logic [39:0] gzdLLzicase67426;
  logic [44:0] callResR7;
  logic [44:0] gzdLLzilambda67423;
  logic [44:0] gzdLLzicase67421;
  logic [39:0] gzdLLzilambda62543;
  logic [46:0] gzdLLzicase67544;
  logic [43:0] gzdLLzicase62547;
  logic [43:0] gMainzislsmzuconnecting;
  logic [68:0] gzdLLzilambda67353;
  logic [68:0] gzdLLzicase67350;
  logic [68:0] gzdLLzilambda63152;
  logic [24:0] gzdLLzicase62969;
  logic [43:0] gzdLLzilambda66854;
  logic [43:0] gzdLLzicase66851;
  logic [43:0] gzdLLzilambda63149;
  logic [68:0] gzdLLzilambda66847;
  logic [68:0] gzdLLzicase66844;
  logic [68:0] gzdLLzilambda63146;
  logic [24:0] gMainzirxzuerrorzusyncR1;
  logic [0:0] callResR8;
  logic [24:0] gMainzirxzuerrorzusyncR2;
  logic [0:0] callResR9;
  logic [69:0] gzdLLzicase66838;
  logic [68:0] gzdLLzicase63139;
  logic [24:0] gMainzilinkzudisablezuzz1R1;
  logic [0:0] callResR10;
  logic [24:0] gMainzilinkzudisablezuzz1R2;
  logic [0:0] callResR11;
  logic [44:0] gzdLLzicase66501;
  logic [43:0] gzdLLzicase63135;
  logic [18:0] gMainziizuafterzu12p8zuus;
  logic [0:0] callResR12;
  logic [18:0] gMainziizuafterzu12p8zuusR1;
  logic [0:0] callResR13;
  logic [44:0] gzdLLzicase66491;
  logic [43:0] gzdLLzicase63132;
  logic [18:0] gMainzigotzunzucharzusync;
  logic [0:0] callResR14;
  logic [18:0] gMainzigotzutimezucodezusync;
  logic [0:0] callResR15;
  logic [1:0] gReWireziPreludezizbzbR2;
  logic [0:0] callResR16;
  logic [18:0] gMainzigotzunzucharzusyncR1;
  logic [0:0] callResR17;
  logic [18:0] gMainzigotzutimezucodezusyncR1;
  logic [0:0] callResR18;
  logic [1:0] gReWireziPreludezizbzbR3;
  logic [0:0] callResR19;
  logic [44:0] gzdLLzicase66481;
  logic [43:0] gzdLLzicase63129;
  logic [18:0] gMainzigotzufctzusync;
  logic [0:0] callResR20;
  logic [18:0] gMainzigotzufctzusyncR1;
  logic [0:0] callResR21;
  logic [25:0] gzdLLzicase66471;
  logic [24:0] gzdLLzicase63126;
  logic [49:0] gzdLLzilambda66464;
  logic [49:0] gzdLLzilambda63125;
  logic [24:0] gzdLLzicase63123;
  logic [24:0] callResR22;
  logic [25:0] gzdLLzicase66473;
  logic [24:0] gzdLLzicase63127;
  logic [49:0] gzdLLzilambda66469;
  logic [49:0] gzdLLzilambda63099;
  logic [24:0] gzdLLzicase63097;
  logic [25:0] gzdLLzicase66483;
  logic [24:0] gzdLLzicase63130;
  logic [49:0] gzdLLzilambda66478;
  logic [49:0] gzdLLzilambda63073;
  logic [24:0] gzdLLzicase63071;
  logic [24:0] callResR23;
  logic [25:0] gzdLLzicase66493;
  logic [24:0] gzdLLzicase63133;
  logic [49:0] gzdLLzilambda66488;
  logic [49:0] gzdLLzilambda63047;
  logic [24:0] gzdLLzicase62993R1;
  logic [24:0] callResR24;
  logic [25:0] gzdLLzicase66503;
  logic [24:0] gzdLLzicase63136;
  logic [49:0] gzdLLzilambda66498;
  logic [49:0] gzdLLzilambda63021;
  logic [24:0] gzdLLzicase62993R2;
  logic [24:0] callResR25;
  logic [25:0] gzdLLzicase66840;
  logic [24:0] gzdLLzicase63140;
  logic [49:0] gzdLLzilambda66508;
  logic [49:0] gzdLLzilambda62995;
  logic [24:0] gzdLLzicase62993R3;
  logic [24:0] callResR26;
  logic [43:0] gzdLLzilambda66834;
  logic [43:0] gzdLLzicase66831R1;
  logic [39:0] callResR27;
  logic [39:0] gzdLLzilambda67438;
  logic [39:0] gzdLLzicase67426R1;
  logic [44:0] callResR28;
  logic [44:0] gzdLLzilambda67433;
  logic [44:0] gzdLLzicase67431;
  logic [39:0] gzdLLzilambda62539;
  logic [46:0] gzdLLzicase67547;
  logic [43:0] gzdLLzicase62549;
  logic [43:0] gMainzislsmzustarted;
  logic [68:0] gzdLLzilambda67413;
  logic [68:0] gzdLLzicase67410;
  logic [68:0] gzdLLzilambda63999;
  logic [24:0] gzdLLzicase63843;
  logic [43:0] gzdLLzilambda67117;
  logic [43:0] gzdLLzicase67114;
  logic [43:0] gzdLLzilambda63996;
  logic [68:0] gzdLLzilambda67110;
  logic [68:0] gzdLLzicase67107;
  logic [68:0] gzdLLzilambda63993;
  logic [24:0] gMainzirxzuerrorzusyncR3;
  logic [0:0] callResR29;
  logic [24:0] gMainzilinkzudisablezuzz1R3;
  logic [0:0] callResR30;
  logic [1:0] gReWireziPreludezizbzbR4;
  logic [0:0] callResR31;
  logic [24:0] gMainzirxzuerrorzusyncR4;
  logic [0:0] callResR32;
  logic [24:0] gMainzilinkzudisablezuzz1R4;
  logic [0:0] callResR33;
  logic [1:0] gReWireziPreludezizbzbR5;
  logic [0:0] callResR34;
  logic [69:0] gzdLLzicase67101;
  logic [68:0] gzdLLzicase63986;
  logic [18:0] gMainzigotzufctzusyncR2;
  logic [0:0] callResR35;
  logic [18:0] gMainzigotzunzucharzusyncR2;
  logic [0:0] callResR36;
  logic [18:0] gMainzigotzutimezucodezusyncR2;
  logic [0:0] callResR37;
  logic [1:0] gReWireziPreludezizbzbR6;
  logic [0:0] callResR38;
  logic [1:0] gReWireziPreludezizbzbR7;
  logic [0:0] callResR39;
  logic [18:0] gMainzigotzufctzusyncR3;
  logic [0:0] callResR40;
  logic [18:0] gMainzigotzunzucharzusyncR3;
  logic [0:0] callResR41;
  logic [18:0] gMainzigotzutimezucodezusyncR3;
  logic [0:0] callResR42;
  logic [1:0] gReWireziPreludezizbzbR8;
  logic [0:0] callResR43;
  logic [1:0] gReWireziPreludezizbzbR9;
  logic [0:0] callResR44;
  logic [69:0] gzdLLzicase66639;
  logic [68:0] gzdLLzicase63982;
  logic [18:0] gMainziizuafterzu12p8zuusR2;
  logic [0:0] callResR45;
  logic [18:0] gMainziizuafterzu12p8zuusR3;
  logic [0:0] callResR46;
  logic [69:0] gzdLLzicase66628;
  logic [68:0] gzdLLzicase63978;
  logic [18:0] gMainzigotzunullzusync;
  logic [0:0] callResR47;
  logic [24:0] gMainzigotzunullzusynczureg;
  logic [0:0] callResR48;
  logic [1:0] gReWireziPreludezizbzbR10;
  logic [0:0] callResR49;
  logic [18:0] gMainzigotzunullzusyncR1;
  logic [0:0] callResR50;
  logic [24:0] gMainzigotzunullzusynczuregR1;
  logic [0:0] callResR51;
  logic [1:0] gReWireziPreludezizbzbR11;
  logic [0:0] callResR52;
  logic [25:0] gzdLLzicase66617;
  logic [24:0] gzdLLzicase63974;
  logic [49:0] gzdLLzilambda66610;
  logic [49:0] gzdLLzilambda63973;
  logic [24:0] gzdLLzicase63123R1;
  logic [24:0] callResR53;
  logic [25:0] gzdLLzicase66619;
  logic [24:0] gzdLLzicase63975;
  logic [49:0] gzdLLzilambda66615;
  logic [49:0] gzdLLzilambda63947;
  logic [24:0] gzdLLzicase63945;
  logic [25:0] gzdLLzicase66630;
  logic [24:0] gzdLLzicase63979;
  logic [49:0] gzdLLzilambda66624;
  logic [49:0] gzdLLzilambda63921;
  logic [24:0] gzdLLzicase62993R4;
  logic [24:0] callResR54;
  logic [25:0] gzdLLzicase66641;
  logic [24:0] gzdLLzicase63983;
  logic [49:0] gzdLLzilambda66635;
  logic [49:0] gzdLLzilambda63895;
  logic [24:0] gzdLLzicase63071R1;
  logic [24:0] callResR55;
  logic [25:0] gzdLLzicase67103;
  logic [24:0] gzdLLzicase63987;
  logic [49:0] gzdLLzilambda66646;
  logic [49:0] gzdLLzilambda63869;
  logic [24:0] gzdLLzicase62993R5;
  logic [24:0] callResR56;
  logic [43:0] gzdLLzilambda67097;
  logic [43:0] gzdLLzicase66831R2;
  logic [39:0] callResR57;
  logic [39:0] gzdLLzilambda67448;
  logic [39:0] gzdLLzicase67426R2;
  logic [44:0] callResR58;
  logic [44:0] gzdLLzilambda67443;
  logic [44:0] gzdLLzicase67441;
  logic [39:0] gzdLLzilambda62535;
  logic [46:0] gzdLLzicase67550;
  logic [43:0] gzdLLzicase62551;
  logic [43:0] gMainzislsmzuready;
  logic [68:0] gzdLLzilambda67389;
  logic [68:0] gzdLLzicase67386;
  logic [68:0] gzdLLzilambda63706;
  logic [24:0] gzdLLzicase63521;
  logic [43:0] gzdLLzilambda67010;
  logic [43:0] gzdLLzicase67007;
  logic [43:0] gzdLLzilambda63703;
  logic [18:0] gMainzigotzunullzusyncR2;
  logic [0:0] callResR59;
  logic [18:0] gMainzigotzunullzusyncR3;
  logic [0:0] callResR60;
  logic [25:0] idR1;
  logic [25:0] gzdLLzicase67003;
  logic [24:0] gzdLLzicase63549;
  logic [49:0] gzdLLzilambda66561;
  logic [49:0] gzdLLzilambda63547;
  logic [24:0] gzdLLzicase63392;
  logic [24:0] callResR61;
  logic [43:0] gzdLLzilambda66999;
  logic [43:0] gzdLLzicase66996;
  logic [43:0] gzdLLzilambda63700;
  logic [68:0] gzdLLzilambda66992;
  logic [68:0] gzdLLzicase66989;
  logic [68:0] gzdLLzilambda63697;
  logic [24:0] gMainzirxzuerrorzusyncR5;
  logic [0:0] callResR62;
  logic [24:0] gMainzirxzuerrorzusyncR6;
  logic [0:0] callResR63;
  logic [69:0] gzdLLzicase66983;
  logic [68:0] gzdLLzicase63690;
  logic [18:0] gMainzigotzufctzusyncR4;
  logic [0:0] callResR64;
  logic [18:0] gMainzigotzunzucharzusyncR4;
  logic [0:0] callResR65;
  logic [18:0] gMainzigotzutimezucodezusyncR4;
  logic [0:0] callResR66;
  logic [1:0] gReWireziPreludezizbzbR12;
  logic [0:0] callResR67;
  logic [1:0] gReWireziPreludezizbzbR13;
  logic [0:0] callResR68;
  logic [18:0] gMainzigotzufctzusyncR5;
  logic [0:0] callResR69;
  logic [18:0] gMainzigotzunzucharzusyncR5;
  logic [0:0] callResR70;
  logic [18:0] gMainzigotzutimezucodezusyncR5;
  logic [0:0] callResR71;
  logic [1:0] gReWireziPreludezizbzbR14;
  logic [0:0] callResR72;
  logic [1:0] gReWireziPreludezizbzbR15;
  logic [0:0] callResR73;
  logic [50:0] gzdLLzicase66593;
  logic [49:0] gzdLLzicase63686;
  logic [24:0] gMainziautozustartzuzz1;
  logic [0:0] callResR74;
  logic [24:0] gMainzigotzunullzusynczuregR2;
  logic [0:0] callResR75;
  logic [1:0] gReWireziPreludezizaza;
  logic [0:0] callResR76;
  logic [24:0] gMainziautozustartzuzz1R1;
  logic [0:0] callResR77;
  logic [24:0] gMainzigotzunullzusynczuregR3;
  logic [0:0] callResR78;
  logic [1:0] gReWireziPreludezizazaR1;
  logic [0:0] callResR79;
  logic [50:0] gzdLLzicase66583;
  logic [49:0] gzdLLzicase63683;
  logic [24:0] gMainzilinkzustartzuzz1;
  logic [0:0] callResR80;
  logic [24:0] gMainzilinkzustartzuzz1R1;
  logic [0:0] callResR81;
  logic [25:0] gzdLLzicase66573;
  logic [24:0] gzdLLzicase63680;
  logic [49:0] gzdLLzilambda66566;
  logic [49:0] gzdLLzilambda63679;
  logic [24:0] gzdLLzicase63123R2;
  logic [24:0] callResR82;
  logic [25:0] gzdLLzicase66575;
  logic [24:0] gzdLLzicase63681;
  logic [49:0] gzdLLzilambda66571;
  logic [49:0] gzdLLzilambda63653;
  logic [24:0] gzdLLzicase63625;
  logic [24:0] callResR83;
  logic [25:0] gzdLLzicase66585;
  logic [24:0] gzdLLzicase63684;
  logic [49:0] gzdLLzilambda66580;
  logic [49:0] gzdLLzilambda63627;
  logic [24:0] gzdLLzicase63625R1;
  logic [24:0] callResR84;
  logic [25:0] gzdLLzicase66595;
  logic [24:0] gzdLLzicase63687;
  logic [49:0] gzdLLzilambda66590;
  logic [49:0] gzdLLzilambda63601;
  logic [24:0] gzdLLzicase63071R2;
  logic [24:0] callResR85;
  logic [25:0] gzdLLzicase66985;
  logic [24:0] gzdLLzicase63691;
  logic [49:0] gzdLLzilambda66600;
  logic [49:0] gzdLLzilambda63575;
  logic [24:0] gzdLLzicase62993R6;
  logic [24:0] callResR86;
  logic [43:0] gzdLLzilambda66979;
  logic [43:0] gzdLLzicase66831R3;
  logic [39:0] callResR87;
  logic [39:0] gzdLLzilambda67458;
  logic [39:0] gzdLLzicase67426R3;
  logic [44:0] callResR88;
  logic [44:0] gzdLLzilambda67453;
  logic [44:0] gzdLLzicase67451;
  logic [39:0] gzdLLzilambda62531;
  logic [46:0] gzdLLzicase67553;
  logic [43:0] gzdLLzicase62553;
  logic [43:0] gMainzislsmzuerrorzuwait;
  logic [68:0] gzdLLzilambda67377;
  logic [68:0] gzdLLzicase67374;
  logic [68:0] gzdLLzilambda63497;
  logic [24:0] gzdLLzicase63368;
  logic [43:0] gzdLLzilambda66972;
  logic [43:0] gzdLLzicase66969;
  logic [43:0] gzdLLzilambda63494;
  logic [18:0] gMainzigotzunullzusyncR4;
  logic [0:0] callResR89;
  logic [18:0] gMainzigotzunullzusyncR5;
  logic [0:0] callResR90;
  logic [25:0] idR2;
  logic [25:0] gzdLLzicase66965;
  logic [24:0] gzdLLzicase63396;
  logic [49:0] gzdLLzilambda66532;
  logic [49:0] gzdLLzilambda63394;
  logic [24:0] gzdLLzicase63392R1;
  logic [24:0] callResR91;
  logic [43:0] gzdLLzilambda66961;
  logic [43:0] gzdLLzicase66958;
  logic [43:0] gzdLLzilambda63491;
  logic [68:0] gzdLLzilambda66954;
  logic [68:0] gzdLLzicase66951;
  logic [68:0] gzdLLzilambda63488;
  logic [24:0] gMainzirxzuerrorzusyncR7;
  logic [0:0] callResR92;
  logic [24:0] gMainzirxzuerrorzusyncR8;
  logic [0:0] callResR93;
  logic [44:0] gzdLLzicase66945;
  logic [43:0] gzdLLzicase63481;
  logic [18:0] gMainzigotzufctzusyncR6;
  logic [0:0] callResR94;
  logic [18:0] gMainzigotzunzucharzusyncR6;
  logic [0:0] callResR95;
  logic [18:0] gMainzigotzutimezucodezusyncR6;
  logic [0:0] callResR96;
  logic [1:0] gReWireziPreludezizbzbR16;
  logic [0:0] callResR97;
  logic [1:0] gReWireziPreludezizbzbR17;
  logic [0:0] callResR98;
  logic [18:0] gMainzigotzufctzusyncR7;
  logic [0:0] callResR99;
  logic [18:0] gMainzigotzunzucharzusyncR7;
  logic [0:0] callResR100;
  logic [18:0] gMainzigotzutimezucodezusyncR7;
  logic [0:0] callResR101;
  logic [1:0] gReWireziPreludezizbzbR18;
  logic [0:0] callResR102;
  logic [1:0] gReWireziPreludezizbzbR19;
  logic [0:0] callResR103;
  logic [44:0] gzdLLzicase66549;
  logic [43:0] gzdLLzicase63478;
  logic [18:0] gMainziizuafterzu12p8zuusR4;
  logic [0:0] callResR104;
  logic [18:0] gMainziizuafterzu12p8zuusR5;
  logic [0:0] callResR105;
  logic [25:0] idR3;
  logic [25:0] gzdLLzicase66541;
  logic [24:0] gzdLLzicase63476;
  logic [49:0] gzdLLzilambda66537;
  logic [49:0] gzdLLzilambda63474;
  logic [24:0] gzdLLzicase63472;
  logic [25:0] gzdLLzicase66551;
  logic [24:0] gzdLLzicase63479;
  logic [49:0] gzdLLzilambda66546;
  logic [49:0] gzdLLzilambda63448;
  logic [24:0] gzdLLzicase63071R3;
  logic [24:0] callResR106;
  logic [25:0] gzdLLzicase66947;
  logic [24:0] gzdLLzicase63482;
  logic [49:0] gzdLLzilambda66556;
  logic [49:0] gzdLLzilambda63422;
  logic [24:0] gzdLLzicase62993R7;
  logic [24:0] callResR107;
  logic [43:0] gzdLLzilambda66942;
  logic [43:0] gzdLLzicase66831R4;
  logic [39:0] callResR108;
  logic [39:0] gzdLLzilambda67468;
  logic [39:0] gzdLLzicase67426R4;
  logic [44:0] callResR109;
  logic [44:0] gzdLLzilambda67463;
  logic [44:0] gzdLLzicase67461;
  logic [39:0] gzdLLzilambda62527;
  logic [46:0] gzdLLzicase67556;
  logic [43:0] gzdLLzicase62555;
  logic [43:0] gMainzislsmzuerrorzureset;
  logic [68:0] gzdLLzilambda67365;
  logic [68:0] gzdLLzicase67362;
  logic [68:0] gzdLLzilambda63344;
  logic [24:0] gzdLLzicase63176;
  logic [43:0] gzdLLzilambda66935;
  logic [43:0] gzdLLzicase66932;
  logic [43:0] gzdLLzilambda63341;
  logic [68:0] gzdLLzilambda66928;
  logic [68:0] gzdLLzicase66925;
  logic [68:0] gzdLLzilambda63338;
  logic [93:0] gzdLLzilambda66921;
  logic [93:0] gzdLLzicase66917;
  logic [93:0] gzdLLzilambda63335;
  logic [49:0] gzdLLzicase63201;
  logic [24:0] gMainzisendzutimezucodeR1;
  logic [0:0] callResR110;
  logic [0:0] litR2;
  logic [43:0] gzdLLzilambda66912;
  logic [43:0] gzdLLzicase66909;
  logic [43:0] gzdLLzilambda63331;
  logic [68:0] gzdLLzilambda66905;
  logic [68:0] gzdLLzicase66902;
  logic [68:0] gzdLLzilambda63328;
  logic [24:0] gMainzififozuavailablezuzz1;
  logic [0:0] callResR111;
  logic [24:0] gMainzififozuavailablezuzz1R1;
  logic [0:0] callResR112;
  logic [25:0] idR4;
  logic [25:0] gzdLLzicase66898;
  logic [24:0] gzdLLzicase63229;
  logic [49:0] gzdLLzilambda66513;
  logic [49:0] gzdLLzilambda63227;
  logic [24:0] gzdLLzicase63225;
  logic [43:0] gzdLLzilambda66894;
  logic [43:0] gzdLLzicase66891;
  logic [43:0] gzdLLzilambda63325;
  logic [68:0] gzdLLzilambda66887;
  logic [68:0] gzdLLzicase66884;
  logic [68:0] gzdLLzilambda63322;
  logic [24:0] gzdLLzicase63253;
  logic [43:0] gzdLLzilambda66880;
  logic [43:0] gzdLLzicase66877;
  logic [43:0] gzdLLzilambda63319;
  logic [68:0] gzdLLzilambda66873;
  logic [68:0] gzdLLzicase66870;
  logic [68:0] gzdLLzilambda63316;
  logic [24:0] gMainzirxzuerrorzusyncR9;
  logic [0:0] callResR113;
  logic [24:0] gMainzirxzuerrorzusyncR10;
  logic [0:0] callResR114;
  logic [44:0] gzdLLzicase66864;
  logic [43:0] gzdLLzicase63309;
  logic [18:0] gMainziizuafterzu6p4zuus;
  logic [0:0] callResR115;
  logic [18:0] gMainziizuafterzu6p4zuusR1;
  logic [0:0] callResR116;
  logic [25:0] idR5;
  logic [25:0] gzdLLzicase66522;
  logic [24:0] gzdLLzicase63307;
  logic [49:0] gzdLLzilambda66518;
  logic [49:0] gzdLLzilambda63305;
  logic [24:0] gzdLLzicase63303;
  logic [25:0] gzdLLzicase66866;
  logic [24:0] gzdLLzicase63310;
  logic [49:0] gzdLLzilambda66527;
  logic [49:0] gzdLLzilambda63279;
  logic [24:0] gzdLLzicase63123R3;
  logic [24:0] callResR117;
  logic [43:0] gzdLLzilambda66861;
  logic [43:0] gzdLLzicase66831R5;
  logic [39:0] callResR118;
  logic [39:0] gzdLLzilambda67478;
  logic [39:0] gzdLLzicase67426R5;
  logic [44:0] callResR119;
  logic [44:0] gzdLLzilambda67473;
  logic [44:0] gzdLLzicase67471;
  logic [39:0] gzdLLzilambda62523;
  assign gMainzidispatch = {arg1, arg0};
  assign gzdLLzilambda67585 = {gMainzidispatch[24:0], gMainzidispatch[24:0]};
  assign gzdLLzilambda62519 = gzdLLzilambda67585[49:0];
  assign gMainzilinkzustate = gzdLLzilambda62519[49:25];
  assign gzdLLzicase62798 = gMainzilinkzustate[24:0];
  assign gzdLLzilambda67580 = {gzdLLzicase62798[2:0], gzdLLzilambda62519[24:0]};
  assign gzdLLzicase67578 = gzdLLzilambda67580[27:0];
  assign gzdLLzilambda67575 = {gMainzidispatch[43:25], {17'h01000, gzdLLzicase67578[27:25], gzdLLzicase67578[24:0]}};
  assign gzdLLzicase67572 = {gzdLLzilambda67575[44:0], gzdLLzilambda67575[63:45]};
  assign gzdLLzilambda62558 = {gzdLLzicase67572[18:0], gzdLLzicase67572[46:44], gzdLLzicase67572[43:19]};
  assign gzdLLzicase67541 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62545 = {gzdLLzicase67541[43:25], gzdLLzicase67541[24:0]};
  assign gMainzislsmzurun = {gzdLLzicase62545[43:25], gzdLLzicase62545[24:0]};
  assign gzdLLzilambda67401 = {gMainzislsmzurun[43:25], gMainzislsmzurun[24:0], gMainzislsmzurun[24:0]};
  assign gzdLLzicase67398 = {gzdLLzilambda67401[49:0], gzdLLzilambda67401[68:50]};
  assign gzdLLzilambda63819 = {gzdLLzicase67398[18:0], gzdLLzicase67398[68:44], gzdLLzicase67398[43:19]};
  assign gzdLLzicase63730 = gzdLLzilambda63819[49:25];
  assign gzdLLzilambda67090 = {gzdLLzilambda63819[68:50], {2'h3, gzdLLzicase63730[22], gzdLLzicase63730[21], gzdLLzicase63730[20], 5'h1f, gzdLLzicase63730[14], gzdLLzicase63730[13], gzdLLzicase63730[12], gzdLLzicase63730[11], gzdLLzicase63730[10], gzdLLzicase63730[9], gzdLLzicase63730[8], gzdLLzicase63730[7], gzdLLzicase63730[6], gzdLLzicase63730[5], gzdLLzicase63730[4], gzdLLzicase63730[3], gzdLLzicase63730[2:0]}};
  assign gzdLLzicase67087 = {gzdLLzilambda67090[24:0], gzdLLzilambda67090[43:25]};
  assign gzdLLzilambda63816 = {gzdLLzicase67087[18:0], gzdLLzicase67087[43:19]};
  assign gzdLLzilambda67083 = {gzdLLzilambda63816[43:25], gzdLLzilambda63816[24:0], gzdLLzilambda63816[24:0]};
  assign gzdLLzicase67080 = {gzdLLzilambda67083[49:0], gzdLLzilambda67083[68:50]};
  assign gzdLLzilambda63813 = {gzdLLzicase67080[18:0], gzdLLzicase67080[68:44], gzdLLzicase67080[43:19]};
  assign gMainzisendzutimezucode = gzdLLzilambda63813[49:25];
  Mainzisendzutimezucode  Mainzisendzutimezucode (gMainzisendzutimezucode[24:0], callRes);
  assign gzdLLzilambda67076 = {gzdLLzilambda63813[68:50], callRes, gzdLLzilambda63813[24:0]};
  assign gzdLLzicase67073 = {gzdLLzilambda67076[25:0], gzdLLzilambda67076[44:26]};
  assign gzdLLzilambda63810 = {gzdLLzicase67073[18:0], gzdLLzicase67073[44], gzdLLzicase67073[43:19]};
  assign gzdLLzilambda67069 = {gzdLLzilambda63810[25], gzdLLzilambda63810[44:26], gzdLLzilambda63810[24:0], gzdLLzilambda63810[24:0]};
  assign gzdLLzicase67065 = {gzdLLzilambda67069[49:0], gzdLLzilambda67069[69], gzdLLzilambda67069[68:50]};
  assign gzdLLzilambda63807 = {gzdLLzicase67065[19], gzdLLzicase67065[18:0], gzdLLzicase67065[69:45], gzdLLzicase67065[44:20]};
  assign gzdLLzicase63755 = {gzdLLzilambda63807[49:25], gzdLLzilambda63807[69]};
  assign gReWireziPreludezinot = gzdLLzicase63755[0];
  assign lit = gReWireziPreludezinot[0];
  assign litR1 = (lit[0] == 1'h1) ? 1'h0 : 1'h1;
  assign gzdLLzilambda67060 = {gzdLLzilambda63807[68:50], {gzdLLzicase63755[25], gzdLLzicase63755[24], gzdLLzicase63755[23], gzdLLzicase63755[22], gzdLLzicase63755[21], gzdLLzicase63755[20], gzdLLzicase63755[19], gzdLLzicase63755[18], gzdLLzicase63755[17], gzdLLzicase63755[16], gzdLLzicase63755[15], (litR1[0] == 1'h1) ? 1'h1 : 1'h0, gzdLLzicase63755[13], gzdLLzicase63755[12], gzdLLzicase63755[11], gzdLLzicase63755[10], gzdLLzicase63755[9], gzdLLzicase63755[8], gzdLLzicase63755[7], gzdLLzicase63755[6], gzdLLzicase63755[5], gzdLLzicase63755[4], gzdLLzicase63755[3:1]}};
  assign gzdLLzicase67057 = {gzdLLzilambda67060[24:0], gzdLLzilambda67060[43:25]};
  assign gzdLLzilambda63803 = {gzdLLzicase67057[18:0], gzdLLzicase67057[43:19]};
  assign gzdLLzilambda67053 = {gzdLLzilambda63803[43:25], gzdLLzilambda63803[24:0], gzdLLzilambda63803[24:0]};
  assign gzdLLzicase67050 = {gzdLLzilambda67053[49:0], gzdLLzilambda67053[68:50]};
  assign gzdLLzilambda63800 = {gzdLLzicase67050[18:0], gzdLLzicase67050[68:44], gzdLLzicase67050[43:19]};
  assign gMainzilinkzudisablezuzz1 = gzdLLzilambda63800[49:25];
  Mainzilinkzudisablezuzz1  Mainzilinkzudisablezuzz1 (gMainzilinkzudisablezuzz1[24:0], callResR1);
  assign gzdLLzilambda67046 = {gzdLLzilambda63800[68:50], callResR1, gzdLLzilambda63800[24:0]};
  assign gzdLLzicase67043 = {gzdLLzilambda67046[25:0], gzdLLzilambda67046[44:26]};
  assign gzdLLzilambda63797 = {gzdLLzicase67043[18:0], gzdLLzicase67043[44], gzdLLzicase67043[43:19]};
  assign gzdLLzilambda67039 = {gzdLLzilambda63797[25], gzdLLzilambda63797[44:26], gzdLLzilambda63797[24:0], gzdLLzilambda63797[24:0]};
  assign gzdLLzicase67035 = {gzdLLzilambda67039[49:0], gzdLLzilambda67039[69], gzdLLzilambda67039[68:50]};
  assign gzdLLzilambda63794 = {gzdLLzicase67035[19], gzdLLzicase67035[18:0], gzdLLzicase67035[69:45], gzdLLzicase67035[44:20]};
  assign gMainzirxzuerrorzusync = gzdLLzilambda63794[49:25];
  Mainzirxzuerrorzusync  Mainzirxzuerrorzusync (gMainzirxzuerrorzusync[24:0], callResR2);
  assign gzdLLzilambda67030 = {gzdLLzilambda63794[69], gzdLLzilambda63794[68:50], callResR2, gzdLLzilambda63794[24:0]};
  assign gzdLLzicase67026 = {gzdLLzilambda67030[25:0], gzdLLzilambda67030[45], gzdLLzilambda67030[44:26]};
  assign gzdLLzilambda63790 = {gzdLLzicase67026[19], gzdLLzicase67026[18:0], gzdLLzicase67026[45], gzdLLzicase67026[44:20]};
  assign gReWireziPreludezizbzb = {gzdLLzilambda63790[45], gzdLLzilambda63790[25]};
  ReWireziPreludezizbzb  ReWireziPreludezizbzb (gReWireziPreludezizbzb[1], gReWireziPreludezizbzb[0], callResR3);
  assign gReWireziPreludezizbzbR1 = {gzdLLzilambda63790[45], gzdLLzilambda63790[25]};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR1 (gReWireziPreludezizbzbR1[1], gReWireziPreludezizbzbR1[0], callResR4);
  assign id = {callResR4, gzdLLzilambda63790[24:0]};
  assign gzdLLzicase67021 = {callResR3, gzdLLzilambda63790[24:0]};
  assign gzdLLzicase63783 = gzdLLzicase67021[24:0];
  assign gzdLLzilambda66605 = {gzdLLzicase63783[24:0], gzdLLzicase63783[24:0]};
  assign gzdLLzilambda63781 = gzdLLzilambda66605[49:0];
  assign gzdLLzicase62993 = gzdLLzilambda63781[49:25];
  zdLLzicase62993  zdLLzicase62993 (gzdLLzicase62993[24], gzdLLzicase62993[23], gzdLLzicase62993[22], gzdLLzicase62993[21], gzdLLzicase62993[20], gzdLLzicase62993[19], gzdLLzicase62993[18], gzdLLzicase62993[17], gzdLLzicase62993[16], gzdLLzicase62993[15], gzdLLzicase62993[14], gzdLLzicase62993[13], gzdLLzicase62993[12], gzdLLzicase62993[11], gzdLLzicase62993[10], gzdLLzicase62993[9], gzdLLzicase62993[8], gzdLLzicase62993[7], gzdLLzicase62993[6], gzdLLzicase62993[5], gzdLLzicase62993[4], gzdLLzicase62993[3], gzdLLzicase62993[2:0], callResR5);
  assign gzdLLzilambda67017 = {gzdLLzilambda63790[44:26], (gzdLLzicase67021[25] == 1'h1) ? callResR5 : id[24:0]};
  assign gzdLLzicase66831 = {gzdLLzilambda67017[24:0], gzdLLzilambda67017[43:25]};
  zdLLzicase66831  zdLLzicase66831 (gzdLLzicase66831[43:19], gzdLLzicase66831[18:0], callResR6);
  assign gzdLLzilambda67428 = callResR6;
  assign gzdLLzicase67426 = gzdLLzilambda67428[39:0];
  zdLLzicase67426  zdLLzicase67426 (gzdLLzicase67426[39:25], gzdLLzicase67426[24:0], callResR7);
  assign gzdLLzilambda67423 = callResR7;
  assign gzdLLzicase67421 = gzdLLzilambda67423[44:0];
  assign gzdLLzilambda62543 = {gzdLLzicase67421[39:25], gzdLLzicase67421[24:0]};
  assign gzdLLzicase67544 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62547 = {gzdLLzicase67544[43:25], gzdLLzicase67544[24:0]};
  assign gMainzislsmzuconnecting = {gzdLLzicase62547[43:25], gzdLLzicase62547[24:0]};
  assign gzdLLzilambda67353 = {gMainzislsmzuconnecting[43:25], gMainzislsmzuconnecting[24:0], gMainzislsmzuconnecting[24:0]};
  assign gzdLLzicase67350 = {gzdLLzilambda67353[49:0], gzdLLzilambda67353[68:50]};
  assign gzdLLzilambda63152 = {gzdLLzicase67350[18:0], gzdLLzicase67350[68:44], gzdLLzicase67350[43:19]};
  assign gzdLLzicase62969 = gzdLLzilambda63152[49:25];
  assign gzdLLzilambda66854 = {gzdLLzilambda63152[68:50], {2'h3, gzdLLzicase62969[22], gzdLLzicase62969[21], 3'h3, gzdLLzicase62969[17], gzdLLzicase62969[16], gzdLLzicase62969[15], gzdLLzicase62969[14], gzdLLzicase62969[13], gzdLLzicase62969[12], gzdLLzicase62969[11], gzdLLzicase62969[10], gzdLLzicase62969[9], gzdLLzicase62969[8], gzdLLzicase62969[7], gzdLLzicase62969[6], gzdLLzicase62969[5], gzdLLzicase62969[4], gzdLLzicase62969[3], gzdLLzicase62969[2:0]}};
  assign gzdLLzicase66851 = {gzdLLzilambda66854[24:0], gzdLLzilambda66854[43:25]};
  assign gzdLLzilambda63149 = {gzdLLzicase66851[18:0], gzdLLzicase66851[43:19]};
  assign gzdLLzilambda66847 = {gzdLLzilambda63149[43:25], gzdLLzilambda63149[24:0], gzdLLzilambda63149[24:0]};
  assign gzdLLzicase66844 = {gzdLLzilambda66847[49:0], gzdLLzilambda66847[68:50]};
  assign gzdLLzilambda63146 = {gzdLLzicase66844[18:0], gzdLLzicase66844[68:44], gzdLLzicase66844[43:19]};
  assign gMainzirxzuerrorzusyncR1 = gzdLLzilambda63146[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR1 (gMainzirxzuerrorzusyncR1[24:0], callResR8);
  assign gMainzirxzuerrorzusyncR2 = gzdLLzilambda63146[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR2 (gMainzirxzuerrorzusyncR2[24:0], callResR9);
  assign gzdLLzicase66838 = {callResR9, gzdLLzilambda63146[49:25], gzdLLzilambda63146[68:50], gzdLLzilambda63146[24:0]};
  assign gzdLLzicase63139 = {gzdLLzicase66838[68:44], gzdLLzicase66838[43:25], gzdLLzicase66838[24:0]};
  assign gMainzilinkzudisablezuzz1R1 = gzdLLzicase63139[68:44];
  Mainzilinkzudisablezuzz1  Mainzilinkzudisablezuzz1R1 (gMainzilinkzudisablezuzz1R1[24:0], callResR10);
  assign gMainzilinkzudisablezuzz1R2 = gzdLLzicase63139[68:44];
  Mainzilinkzudisablezuzz1  Mainzilinkzudisablezuzz1R2 (gMainzilinkzudisablezuzz1R2[24:0], callResR11);
  assign gzdLLzicase66501 = {callResR11, gzdLLzicase63139[43:25], gzdLLzicase63139[24:0]};
  assign gzdLLzicase63135 = {gzdLLzicase66501[43:25], gzdLLzicase66501[24:0]};
  assign gMainziizuafterzu12p8zuus = gzdLLzicase63135[43:25];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuus (gMainziizuafterzu12p8zuus[18:0], callResR12);
  assign gMainziizuafterzu12p8zuusR1 = gzdLLzicase63135[43:25];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuusR1 (gMainziizuafterzu12p8zuusR1[18:0], callResR13);
  assign gzdLLzicase66491 = {callResR13, gzdLLzicase63135[43:25], gzdLLzicase63135[24:0]};
  assign gzdLLzicase63132 = {gzdLLzicase66491[43:25], gzdLLzicase66491[24:0]};
  assign gMainzigotzunzucharzusync = gzdLLzicase63132[43:25];
  Mainzigotzunzucharzusync  Mainzigotzunzucharzusync (gMainzigotzunzucharzusync[18:0], callResR14);
  assign gMainzigotzutimezucodezusync = gzdLLzicase63132[43:25];
  Mainzigotzutimezucodezusync  Mainzigotzutimezucodezusync (gMainzigotzutimezucodezusync[18:0], callResR15);
  assign gReWireziPreludezizbzbR2 = {callResR14, callResR15};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR2 (gReWireziPreludezizbzbR2[1], gReWireziPreludezizbzbR2[0], callResR16);
  assign gMainzigotzunzucharzusyncR1 = gzdLLzicase63132[43:25];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR1 (gMainzigotzunzucharzusyncR1[18:0], callResR17);
  assign gMainzigotzutimezucodezusyncR1 = gzdLLzicase63132[43:25];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR1 (gMainzigotzutimezucodezusyncR1[18:0], callResR18);
  assign gReWireziPreludezizbzbR3 = {callResR17, callResR18};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR3 (gReWireziPreludezizbzbR3[1], gReWireziPreludezizbzbR3[0], callResR19);
  assign gzdLLzicase66481 = {callResR19, gzdLLzicase63132[43:25], gzdLLzicase63132[24:0]};
  assign gzdLLzicase63129 = {gzdLLzicase66481[43:25], gzdLLzicase66481[24:0]};
  assign gMainzigotzufctzusync = gzdLLzicase63129[43:25];
  Mainzigotzufctzusync  Mainzigotzufctzusync (gMainzigotzufctzusync[18:0], callResR20);
  assign gMainzigotzufctzusyncR1 = gzdLLzicase63129[43:25];
  Mainzigotzufctzusync  MainzigotzufctzusyncR1 (gMainzigotzufctzusyncR1[18:0], callResR21);
  assign gzdLLzicase66471 = {callResR21, gzdLLzicase63129[24:0]};
  assign gzdLLzicase63126 = gzdLLzicase66471[24:0];
  assign gzdLLzilambda66464 = {gzdLLzicase63126[24:0], gzdLLzicase63126[24:0]};
  assign gzdLLzilambda63125 = gzdLLzilambda66464[49:0];
  assign gzdLLzicase63123 = gzdLLzilambda63125[49:25];
  zdLLzicase63123  zdLLzicase63123 (gzdLLzicase63123[24], gzdLLzicase63123[23], gzdLLzicase63123[22], gzdLLzicase63123[21], gzdLLzicase63123[20], gzdLLzicase63123[19], gzdLLzicase63123[18], gzdLLzicase63123[17], gzdLLzicase63123[16], gzdLLzicase63123[15], gzdLLzicase63123[14], gzdLLzicase63123[13], gzdLLzicase63123[12], gzdLLzicase63123[11], gzdLLzicase63123[10], gzdLLzicase63123[9], gzdLLzicase63123[8], gzdLLzicase63123[7], gzdLLzicase63123[6], gzdLLzicase63123[5], gzdLLzicase63123[4], gzdLLzicase63123[3], gzdLLzicase63123[2:0], callResR22);
  assign gzdLLzicase66473 = {callResR20, gzdLLzicase63129[24:0]};
  assign gzdLLzicase63127 = gzdLLzicase66473[24:0];
  assign gzdLLzilambda66469 = {gzdLLzicase63127[24:0], gzdLLzicase63127[24:0]};
  assign gzdLLzilambda63099 = gzdLLzilambda66469[49:0];
  assign gzdLLzicase63097 = gzdLLzilambda63099[49:25];
  assign gzdLLzicase66483 = {callResR16, gzdLLzicase63132[24:0]};
  assign gzdLLzicase63130 = gzdLLzicase66483[24:0];
  assign gzdLLzilambda66478 = {gzdLLzicase63130[24:0], gzdLLzicase63130[24:0]};
  assign gzdLLzilambda63073 = gzdLLzilambda66478[49:0];
  assign gzdLLzicase63071 = gzdLLzilambda63073[49:25];
  zdLLzicase63071  zdLLzicase63071 (gzdLLzicase63071[24], gzdLLzicase63071[23], gzdLLzicase63071[22], gzdLLzicase63071[21], gzdLLzicase63071[20], gzdLLzicase63071[19], gzdLLzicase63071[18], gzdLLzicase63071[17], gzdLLzicase63071[16], gzdLLzicase63071[15], gzdLLzicase63071[14], gzdLLzicase63071[13], gzdLLzicase63071[12], gzdLLzicase63071[11], gzdLLzicase63071[10], gzdLLzicase63071[9], gzdLLzicase63071[8], gzdLLzicase63071[7], gzdLLzicase63071[6], gzdLLzicase63071[5], gzdLLzicase63071[4], gzdLLzicase63071[3], gzdLLzicase63071[2:0], callResR23);
  assign gzdLLzicase66493 = {callResR12, gzdLLzicase63135[24:0]};
  assign gzdLLzicase63133 = gzdLLzicase66493[24:0];
  assign gzdLLzilambda66488 = {gzdLLzicase63133[24:0], gzdLLzicase63133[24:0]};
  assign gzdLLzilambda63047 = gzdLLzilambda66488[49:0];
  assign gzdLLzicase62993R1 = gzdLLzilambda63047[49:25];
  zdLLzicase62993  zdLLzicase62993R1 (gzdLLzicase62993R1[24], gzdLLzicase62993R1[23], gzdLLzicase62993R1[22], gzdLLzicase62993R1[21], gzdLLzicase62993R1[20], gzdLLzicase62993R1[19], gzdLLzicase62993R1[18], gzdLLzicase62993R1[17], gzdLLzicase62993R1[16], gzdLLzicase62993R1[15], gzdLLzicase62993R1[14], gzdLLzicase62993R1[13], gzdLLzicase62993R1[12], gzdLLzicase62993R1[11], gzdLLzicase62993R1[10], gzdLLzicase62993R1[9], gzdLLzicase62993R1[8], gzdLLzicase62993R1[7], gzdLLzicase62993R1[6], gzdLLzicase62993R1[5], gzdLLzicase62993R1[4], gzdLLzicase62993R1[3], gzdLLzicase62993R1[2:0], callResR24);
  assign gzdLLzicase66503 = {callResR10, gzdLLzicase63139[24:0]};
  assign gzdLLzicase63136 = gzdLLzicase66503[24:0];
  assign gzdLLzilambda66498 = {gzdLLzicase63136[24:0], gzdLLzicase63136[24:0]};
  assign gzdLLzilambda63021 = gzdLLzilambda66498[49:0];
  assign gzdLLzicase62993R2 = gzdLLzilambda63021[49:25];
  zdLLzicase62993  zdLLzicase62993R2 (gzdLLzicase62993R2[24], gzdLLzicase62993R2[23], gzdLLzicase62993R2[22], gzdLLzicase62993R2[21], gzdLLzicase62993R2[20], gzdLLzicase62993R2[19], gzdLLzicase62993R2[18], gzdLLzicase62993R2[17], gzdLLzicase62993R2[16], gzdLLzicase62993R2[15], gzdLLzicase62993R2[14], gzdLLzicase62993R2[13], gzdLLzicase62993R2[12], gzdLLzicase62993R2[11], gzdLLzicase62993R2[10], gzdLLzicase62993R2[9], gzdLLzicase62993R2[8], gzdLLzicase62993R2[7], gzdLLzicase62993R2[6], gzdLLzicase62993R2[5], gzdLLzicase62993R2[4], gzdLLzicase62993R2[3], gzdLLzicase62993R2[2:0], callResR25);
  assign gzdLLzicase66840 = {callResR8, gzdLLzilambda63146[24:0]};
  assign gzdLLzicase63140 = gzdLLzicase66840[24:0];
  assign gzdLLzilambda66508 = {gzdLLzicase63140[24:0], gzdLLzicase63140[24:0]};
  assign gzdLLzilambda62995 = gzdLLzilambda66508[49:0];
  assign gzdLLzicase62993R3 = gzdLLzilambda62995[49:25];
  zdLLzicase62993  zdLLzicase62993R3 (gzdLLzicase62993R3[24], gzdLLzicase62993R3[23], gzdLLzicase62993R3[22], gzdLLzicase62993R3[21], gzdLLzicase62993R3[20], gzdLLzicase62993R3[19], gzdLLzicase62993R3[18], gzdLLzicase62993R3[17], gzdLLzicase62993R3[16], gzdLLzicase62993R3[15], gzdLLzicase62993R3[14], gzdLLzicase62993R3[13], gzdLLzicase62993R3[12], gzdLLzicase62993R3[11], gzdLLzicase62993R3[10], gzdLLzicase62993R3[9], gzdLLzicase62993R3[8], gzdLLzicase62993R3[7], gzdLLzicase62993R3[6], gzdLLzicase62993R3[5], gzdLLzicase62993R3[4], gzdLLzicase62993R3[3], gzdLLzicase62993R3[2:0], callResR26);
  assign gzdLLzilambda66834 = {gzdLLzilambda63146[68:50], (gzdLLzicase66840[25] == 1'h1) ? callResR26 : ((gzdLLzicase66503[25] == 1'h1) ? callResR25 : ((gzdLLzicase66493[25] == 1'h1) ? callResR24 : ((gzdLLzicase66483[25] == 1'h1) ? callResR23 : ((gzdLLzicase66473[25] == 1'h1) ? {gzdLLzicase63097[24], gzdLLzicase63097[23], gzdLLzicase63097[22], gzdLLzicase63097[21], gzdLLzicase63097[20], gzdLLzicase63097[19], gzdLLzicase63097[18], gzdLLzicase63097[17], gzdLLzicase63097[16], gzdLLzicase63097[15], gzdLLzicase63097[14], gzdLLzicase63097[13], gzdLLzicase63097[12], gzdLLzicase63097[11], gzdLLzicase63097[10], gzdLLzicase63097[9], gzdLLzicase63097[8], gzdLLzicase63097[7], gzdLLzicase63097[6], gzdLLzicase63097[5], gzdLLzicase63097[4], gzdLLzicase63097[3], 3'h5} : callResR22))))};
  assign gzdLLzicase66831R1 = {gzdLLzilambda66834[24:0], gzdLLzilambda66834[43:25]};
  zdLLzicase66831  zdLLzicase66831R1 (gzdLLzicase66831R1[43:19], gzdLLzicase66831R1[18:0], callResR27);
  assign gzdLLzilambda67438 = callResR27;
  assign gzdLLzicase67426R1 = gzdLLzilambda67438[39:0];
  zdLLzicase67426  zdLLzicase67426R1 (gzdLLzicase67426R1[39:25], gzdLLzicase67426R1[24:0], callResR28);
  assign gzdLLzilambda67433 = callResR28;
  assign gzdLLzicase67431 = gzdLLzilambda67433[44:0];
  assign gzdLLzilambda62539 = {gzdLLzicase67431[39:25], gzdLLzicase67431[24:0]};
  assign gzdLLzicase67547 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62549 = {gzdLLzicase67547[43:25], gzdLLzicase67547[24:0]};
  assign gMainzislsmzustarted = {gzdLLzicase62549[43:25], gzdLLzicase62549[24:0]};
  assign gzdLLzilambda67413 = {gMainzislsmzustarted[43:25], gMainzislsmzustarted[24:0], gMainzislsmzustarted[24:0]};
  assign gzdLLzicase67410 = {gzdLLzilambda67413[49:0], gzdLLzilambda67413[68:50]};
  assign gzdLLzilambda63999 = {gzdLLzicase67410[18:0], gzdLLzicase67410[68:44], gzdLLzicase67410[43:19]};
  assign gzdLLzicase63843 = gzdLLzilambda63999[49:25];
  assign gzdLLzilambda67117 = {gzdLLzilambda63999[68:50], {2'h3, gzdLLzicase63843[22], gzdLLzicase63843[21], 1'h0, gzdLLzicase63843[19], 1'h1, gzdLLzicase63843[17], gzdLLzicase63843[16], gzdLLzicase63843[15], gzdLLzicase63843[14], gzdLLzicase63843[13], gzdLLzicase63843[12], gzdLLzicase63843[11], gzdLLzicase63843[10], gzdLLzicase63843[9], gzdLLzicase63843[8], gzdLLzicase63843[7], gzdLLzicase63843[6], gzdLLzicase63843[5], gzdLLzicase63843[4], gzdLLzicase63843[3], gzdLLzicase63843[2:0]}};
  assign gzdLLzicase67114 = {gzdLLzilambda67117[24:0], gzdLLzilambda67117[43:25]};
  assign gzdLLzilambda63996 = {gzdLLzicase67114[18:0], gzdLLzicase67114[43:19]};
  assign gzdLLzilambda67110 = {gzdLLzilambda63996[43:25], gzdLLzilambda63996[24:0], gzdLLzilambda63996[24:0]};
  assign gzdLLzicase67107 = {gzdLLzilambda67110[49:0], gzdLLzilambda67110[68:50]};
  assign gzdLLzilambda63993 = {gzdLLzicase67107[18:0], gzdLLzicase67107[68:44], gzdLLzicase67107[43:19]};
  assign gMainzirxzuerrorzusyncR3 = gzdLLzilambda63993[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR3 (gMainzirxzuerrorzusyncR3[24:0], callResR29);
  assign gMainzilinkzudisablezuzz1R3 = gzdLLzilambda63993[49:25];
  Mainzilinkzudisablezuzz1  Mainzilinkzudisablezuzz1R3 (gMainzilinkzudisablezuzz1R3[24:0], callResR30);
  assign gReWireziPreludezizbzbR4 = {callResR29, callResR30};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR4 (gReWireziPreludezizbzbR4[1], gReWireziPreludezizbzbR4[0], callResR31);
  assign gMainzirxzuerrorzusyncR4 = gzdLLzilambda63993[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR4 (gMainzirxzuerrorzusyncR4[24:0], callResR32);
  assign gMainzilinkzudisablezuzz1R4 = gzdLLzilambda63993[49:25];
  Mainzilinkzudisablezuzz1  Mainzilinkzudisablezuzz1R4 (gMainzilinkzudisablezuzz1R4[24:0], callResR33);
  assign gReWireziPreludezizbzbR5 = {callResR32, callResR33};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR5 (gReWireziPreludezizbzbR5[1], gReWireziPreludezizbzbR5[0], callResR34);
  assign gzdLLzicase67101 = {callResR34, gzdLLzilambda63993[68:50], gzdLLzilambda63993[49:25], gzdLLzilambda63993[24:0]};
  assign gzdLLzicase63986 = {gzdLLzicase67101[68:50], gzdLLzicase67101[49:25], gzdLLzicase67101[24:0]};
  assign gMainzigotzufctzusyncR2 = gzdLLzicase63986[68:50];
  Mainzigotzufctzusync  MainzigotzufctzusyncR2 (gMainzigotzufctzusyncR2[18:0], callResR35);
  assign gMainzigotzunzucharzusyncR2 = gzdLLzicase63986[68:50];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR2 (gMainzigotzunzucharzusyncR2[18:0], callResR36);
  assign gMainzigotzutimezucodezusyncR2 = gzdLLzicase63986[68:50];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR2 (gMainzigotzutimezucodezusyncR2[18:0], callResR37);
  assign gReWireziPreludezizbzbR6 = {callResR36, callResR37};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR6 (gReWireziPreludezizbzbR6[1], gReWireziPreludezizbzbR6[0], callResR38);
  assign gReWireziPreludezizbzbR7 = {callResR35, callResR38};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR7 (gReWireziPreludezizbzbR7[1], gReWireziPreludezizbzbR7[0], callResR39);
  assign gMainzigotzufctzusyncR3 = gzdLLzicase63986[68:50];
  Mainzigotzufctzusync  MainzigotzufctzusyncR3 (gMainzigotzufctzusyncR3[18:0], callResR40);
  assign gMainzigotzunzucharzusyncR3 = gzdLLzicase63986[68:50];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR3 (gMainzigotzunzucharzusyncR3[18:0], callResR41);
  assign gMainzigotzutimezucodezusyncR3 = gzdLLzicase63986[68:50];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR3 (gMainzigotzutimezucodezusyncR3[18:0], callResR42);
  assign gReWireziPreludezizbzbR8 = {callResR41, callResR42};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR8 (gReWireziPreludezizbzbR8[1], gReWireziPreludezizbzbR8[0], callResR43);
  assign gReWireziPreludezizbzbR9 = {callResR40, callResR43};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR9 (gReWireziPreludezizbzbR9[1], gReWireziPreludezizbzbR9[0], callResR44);
  assign gzdLLzicase66639 = {callResR44, gzdLLzicase63986[68:50], gzdLLzicase63986[49:25], gzdLLzicase63986[24:0]};
  assign gzdLLzicase63982 = {gzdLLzicase66639[68:50], gzdLLzicase66639[49:25], gzdLLzicase66639[24:0]};
  assign gMainziizuafterzu12p8zuusR2 = gzdLLzicase63982[68:50];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuusR2 (gMainziizuafterzu12p8zuusR2[18:0], callResR45);
  assign gMainziizuafterzu12p8zuusR3 = gzdLLzicase63982[68:50];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuusR3 (gMainziizuafterzu12p8zuusR3[18:0], callResR46);
  assign gzdLLzicase66628 = {callResR46, gzdLLzicase63982[68:50], gzdLLzicase63982[49:25], gzdLLzicase63982[24:0]};
  assign gzdLLzicase63978 = {gzdLLzicase66628[68:50], gzdLLzicase66628[49:25], gzdLLzicase66628[24:0]};
  assign gMainzigotzunullzusync = gzdLLzicase63978[68:50];
  Mainzigotzunullzusync  Mainzigotzunullzusync (gMainzigotzunullzusync[18:0], callResR47);
  assign gMainzigotzunullzusynczureg = gzdLLzicase63978[49:25];
  Mainzigotzunullzusynczureg  Mainzigotzunullzusynczureg (gMainzigotzunullzusynczureg[24:0], callResR48);
  assign gReWireziPreludezizbzbR10 = {callResR47, callResR48};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR10 (gReWireziPreludezizbzbR10[1], gReWireziPreludezizbzbR10[0], callResR49);
  assign gMainzigotzunullzusyncR1 = gzdLLzicase63978[68:50];
  Mainzigotzunullzusync  MainzigotzunullzusyncR1 (gMainzigotzunullzusyncR1[18:0], callResR50);
  assign gMainzigotzunullzusynczuregR1 = gzdLLzicase63978[49:25];
  Mainzigotzunullzusynczureg  MainzigotzunullzusynczuregR1 (gMainzigotzunullzusynczuregR1[24:0], callResR51);
  assign gReWireziPreludezizbzbR11 = {callResR50, callResR51};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR11 (gReWireziPreludezizbzbR11[1], gReWireziPreludezizbzbR11[0], callResR52);
  assign gzdLLzicase66617 = {callResR52, gzdLLzicase63978[24:0]};
  assign gzdLLzicase63974 = gzdLLzicase66617[24:0];
  assign gzdLLzilambda66610 = {gzdLLzicase63974[24:0], gzdLLzicase63974[24:0]};
  assign gzdLLzilambda63973 = gzdLLzilambda66610[49:0];
  assign gzdLLzicase63123R1 = gzdLLzilambda63973[49:25];
  zdLLzicase63123  zdLLzicase63123R1 (gzdLLzicase63123R1[24], gzdLLzicase63123R1[23], gzdLLzicase63123R1[22], gzdLLzicase63123R1[21], gzdLLzicase63123R1[20], gzdLLzicase63123R1[19], gzdLLzicase63123R1[18], gzdLLzicase63123R1[17], gzdLLzicase63123R1[16], gzdLLzicase63123R1[15], gzdLLzicase63123R1[14], gzdLLzicase63123R1[13], gzdLLzicase63123R1[12], gzdLLzicase63123R1[11], gzdLLzicase63123R1[10], gzdLLzicase63123R1[9], gzdLLzicase63123R1[8], gzdLLzicase63123R1[7], gzdLLzicase63123R1[6], gzdLLzicase63123R1[5], gzdLLzicase63123R1[4], gzdLLzicase63123R1[3], gzdLLzicase63123R1[2:0], callResR53);
  assign gzdLLzicase66619 = {callResR49, gzdLLzicase63978[24:0]};
  assign gzdLLzicase63975 = gzdLLzicase66619[24:0];
  assign gzdLLzilambda66615 = {gzdLLzicase63975[24:0], gzdLLzicase63975[24:0]};
  assign gzdLLzilambda63947 = gzdLLzilambda66615[49:0];
  assign gzdLLzicase63945 = gzdLLzilambda63947[49:25];
  assign gzdLLzicase66630 = {callResR45, gzdLLzicase63982[24:0]};
  assign gzdLLzicase63979 = gzdLLzicase66630[24:0];
  assign gzdLLzilambda66624 = {gzdLLzicase63979[24:0], gzdLLzicase63979[24:0]};
  assign gzdLLzilambda63921 = gzdLLzilambda66624[49:0];
  assign gzdLLzicase62993R4 = gzdLLzilambda63921[49:25];
  zdLLzicase62993  zdLLzicase62993R4 (gzdLLzicase62993R4[24], gzdLLzicase62993R4[23], gzdLLzicase62993R4[22], gzdLLzicase62993R4[21], gzdLLzicase62993R4[20], gzdLLzicase62993R4[19], gzdLLzicase62993R4[18], gzdLLzicase62993R4[17], gzdLLzicase62993R4[16], gzdLLzicase62993R4[15], gzdLLzicase62993R4[14], gzdLLzicase62993R4[13], gzdLLzicase62993R4[12], gzdLLzicase62993R4[11], gzdLLzicase62993R4[10], gzdLLzicase62993R4[9], gzdLLzicase62993R4[8], gzdLLzicase62993R4[7], gzdLLzicase62993R4[6], gzdLLzicase62993R4[5], gzdLLzicase62993R4[4], gzdLLzicase62993R4[3], gzdLLzicase62993R4[2:0], callResR54);
  assign gzdLLzicase66641 = {callResR39, gzdLLzicase63986[24:0]};
  assign gzdLLzicase63983 = gzdLLzicase66641[24:0];
  assign gzdLLzilambda66635 = {gzdLLzicase63983[24:0], gzdLLzicase63983[24:0]};
  assign gzdLLzilambda63895 = gzdLLzilambda66635[49:0];
  assign gzdLLzicase63071R1 = gzdLLzilambda63895[49:25];
  zdLLzicase63071  zdLLzicase63071R1 (gzdLLzicase63071R1[24], gzdLLzicase63071R1[23], gzdLLzicase63071R1[22], gzdLLzicase63071R1[21], gzdLLzicase63071R1[20], gzdLLzicase63071R1[19], gzdLLzicase63071R1[18], gzdLLzicase63071R1[17], gzdLLzicase63071R1[16], gzdLLzicase63071R1[15], gzdLLzicase63071R1[14], gzdLLzicase63071R1[13], gzdLLzicase63071R1[12], gzdLLzicase63071R1[11], gzdLLzicase63071R1[10], gzdLLzicase63071R1[9], gzdLLzicase63071R1[8], gzdLLzicase63071R1[7], gzdLLzicase63071R1[6], gzdLLzicase63071R1[5], gzdLLzicase63071R1[4], gzdLLzicase63071R1[3], gzdLLzicase63071R1[2:0], callResR55);
  assign gzdLLzicase67103 = {callResR31, gzdLLzilambda63993[24:0]};
  assign gzdLLzicase63987 = gzdLLzicase67103[24:0];
  assign gzdLLzilambda66646 = {gzdLLzicase63987[24:0], gzdLLzicase63987[24:0]};
  assign gzdLLzilambda63869 = gzdLLzilambda66646[49:0];
  assign gzdLLzicase62993R5 = gzdLLzilambda63869[49:25];
  zdLLzicase62993  zdLLzicase62993R5 (gzdLLzicase62993R5[24], gzdLLzicase62993R5[23], gzdLLzicase62993R5[22], gzdLLzicase62993R5[21], gzdLLzicase62993R5[20], gzdLLzicase62993R5[19], gzdLLzicase62993R5[18], gzdLLzicase62993R5[17], gzdLLzicase62993R5[16], gzdLLzicase62993R5[15], gzdLLzicase62993R5[14], gzdLLzicase62993R5[13], gzdLLzicase62993R5[12], gzdLLzicase62993R5[11], gzdLLzicase62993R5[10], gzdLLzicase62993R5[9], gzdLLzicase62993R5[8], gzdLLzicase62993R5[7], gzdLLzicase62993R5[6], gzdLLzicase62993R5[5], gzdLLzicase62993R5[4], gzdLLzicase62993R5[3], gzdLLzicase62993R5[2:0], callResR56);
  assign gzdLLzilambda67097 = {gzdLLzilambda63993[68:50], (gzdLLzicase67103[25] == 1'h1) ? callResR56 : ((gzdLLzicase66641[25] == 1'h1) ? callResR55 : ((gzdLLzicase66630[25] == 1'h1) ? callResR54 : ((gzdLLzicase66619[25] == 1'h1) ? {gzdLLzicase63945[24], gzdLLzicase63945[23], gzdLLzicase63945[22], gzdLLzicase63945[21], 1'h1, gzdLLzicase63945[19], gzdLLzicase63945[18], gzdLLzicase63945[17], gzdLLzicase63945[16], gzdLLzicase63945[15], gzdLLzicase63945[14], gzdLLzicase63945[13], gzdLLzicase63945[12], gzdLLzicase63945[11], gzdLLzicase63945[10], gzdLLzicase63945[9], gzdLLzicase63945[8], gzdLLzicase63945[7], gzdLLzicase63945[6], gzdLLzicase63945[5], gzdLLzicase63945[4], gzdLLzicase63945[3], 3'h4} : callResR53)))};
  assign gzdLLzicase66831R2 = {gzdLLzilambda67097[24:0], gzdLLzilambda67097[43:25]};
  zdLLzicase66831  zdLLzicase66831R2 (gzdLLzicase66831R2[43:19], gzdLLzicase66831R2[18:0], callResR57);
  assign gzdLLzilambda67448 = callResR57;
  assign gzdLLzicase67426R2 = gzdLLzilambda67448[39:0];
  zdLLzicase67426  zdLLzicase67426R2 (gzdLLzicase67426R2[39:25], gzdLLzicase67426R2[24:0], callResR58);
  assign gzdLLzilambda67443 = callResR58;
  assign gzdLLzicase67441 = gzdLLzilambda67443[44:0];
  assign gzdLLzilambda62535 = {gzdLLzicase67441[39:25], gzdLLzicase67441[24:0]};
  assign gzdLLzicase67550 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62551 = {gzdLLzicase67550[43:25], gzdLLzicase67550[24:0]};
  assign gMainzislsmzuready = {gzdLLzicase62551[43:25], gzdLLzicase62551[24:0]};
  assign gzdLLzilambda67389 = {gMainzislsmzuready[43:25], gMainzislsmzuready[24:0], gMainzislsmzuready[24:0]};
  assign gzdLLzicase67386 = {gzdLLzilambda67389[49:0], gzdLLzilambda67389[68:50]};
  assign gzdLLzilambda63706 = {gzdLLzicase67386[18:0], gzdLLzicase67386[68:44], gzdLLzicase67386[43:19]};
  assign gzdLLzicase63521 = gzdLLzilambda63706[49:25];
  assign gzdLLzilambda67010 = {gzdLLzilambda63706[68:50], {2'h2, gzdLLzicase63521[22], gzdLLzicase63521[21], gzdLLzicase63521[20], gzdLLzicase63521[19], gzdLLzicase63521[18], gzdLLzicase63521[17], gzdLLzicase63521[16], gzdLLzicase63521[15], gzdLLzicase63521[14], gzdLLzicase63521[13], gzdLLzicase63521[12], gzdLLzicase63521[11], gzdLLzicase63521[10], gzdLLzicase63521[9], gzdLLzicase63521[8], gzdLLzicase63521[7], gzdLLzicase63521[6], gzdLLzicase63521[5], gzdLLzicase63521[4], gzdLLzicase63521[3], gzdLLzicase63521[2:0]}};
  assign gzdLLzicase67007 = {gzdLLzilambda67010[24:0], gzdLLzilambda67010[43:25]};
  assign gzdLLzilambda63703 = {gzdLLzicase67007[18:0], gzdLLzicase67007[43:19]};
  assign gMainzigotzunullzusyncR2 = gzdLLzilambda63703[43:25];
  Mainzigotzunullzusync  MainzigotzunullzusyncR2 (gMainzigotzunullzusyncR2[18:0], callResR59);
  assign gMainzigotzunullzusyncR3 = gzdLLzilambda63703[43:25];
  Mainzigotzunullzusync  MainzigotzunullzusyncR3 (gMainzigotzunullzusyncR3[18:0], callResR60);
  assign idR1 = {callResR60, gzdLLzilambda63703[24:0]};
  assign gzdLLzicase67003 = {callResR59, gzdLLzilambda63703[24:0]};
  assign gzdLLzicase63549 = gzdLLzicase67003[24:0];
  assign gzdLLzilambda66561 = {gzdLLzicase63549[24:0], gzdLLzicase63549[24:0]};
  assign gzdLLzilambda63547 = gzdLLzilambda66561[49:0];
  assign gzdLLzicase63392 = gzdLLzilambda63547[49:25];
  zdLLzicase63392  zdLLzicase63392 (gzdLLzicase63392[24], gzdLLzicase63392[23], gzdLLzicase63392[22], gzdLLzicase63392[21], gzdLLzicase63392[20], gzdLLzicase63392[19], gzdLLzicase63392[18], gzdLLzicase63392[17], gzdLLzicase63392[16], gzdLLzicase63392[15], gzdLLzicase63392[14], gzdLLzicase63392[13], gzdLLzicase63392[12], gzdLLzicase63392[11], gzdLLzicase63392[10], gzdLLzicase63392[9], gzdLLzicase63392[8], gzdLLzicase63392[7], gzdLLzicase63392[6], gzdLLzicase63392[5], gzdLLzicase63392[4], gzdLLzicase63392[3], gzdLLzicase63392[2:0], callResR61);
  assign gzdLLzilambda66999 = {gzdLLzilambda63703[43:25], (gzdLLzicase67003[25] == 1'h1) ? callResR61 : idR1[24:0]};
  assign gzdLLzicase66996 = {gzdLLzilambda66999[24:0], gzdLLzilambda66999[43:25]};
  assign gzdLLzilambda63700 = {gzdLLzicase66996[18:0], gzdLLzicase66996[43:19]};
  assign gzdLLzilambda66992 = {gzdLLzilambda63700[43:25], gzdLLzilambda63700[24:0], gzdLLzilambda63700[24:0]};
  assign gzdLLzicase66989 = {gzdLLzilambda66992[49:0], gzdLLzilambda66992[68:50]};
  assign gzdLLzilambda63697 = {gzdLLzicase66989[18:0], gzdLLzicase66989[68:44], gzdLLzicase66989[43:19]};
  assign gMainzirxzuerrorzusyncR5 = gzdLLzilambda63697[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR5 (gMainzirxzuerrorzusyncR5[24:0], callResR62);
  assign gMainzirxzuerrorzusyncR6 = gzdLLzilambda63697[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR6 (gMainzirxzuerrorzusyncR6[24:0], callResR63);
  assign gzdLLzicase66983 = {callResR63, gzdLLzilambda63697[68:50], gzdLLzilambda63697[49:25], gzdLLzilambda63697[24:0]};
  assign gzdLLzicase63690 = {gzdLLzicase66983[68:50], gzdLLzicase66983[49:25], gzdLLzicase66983[24:0]};
  assign gMainzigotzufctzusyncR4 = gzdLLzicase63690[68:50];
  Mainzigotzufctzusync  MainzigotzufctzusyncR4 (gMainzigotzufctzusyncR4[18:0], callResR64);
  assign gMainzigotzunzucharzusyncR4 = gzdLLzicase63690[68:50];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR4 (gMainzigotzunzucharzusyncR4[18:0], callResR65);
  assign gMainzigotzutimezucodezusyncR4 = gzdLLzicase63690[68:50];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR4 (gMainzigotzutimezucodezusyncR4[18:0], callResR66);
  assign gReWireziPreludezizbzbR12 = {callResR65, callResR66};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR12 (gReWireziPreludezizbzbR12[1], gReWireziPreludezizbzbR12[0], callResR67);
  assign gReWireziPreludezizbzbR13 = {callResR64, callResR67};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR13 (gReWireziPreludezizbzbR13[1], gReWireziPreludezizbzbR13[0], callResR68);
  assign gMainzigotzufctzusyncR5 = gzdLLzicase63690[68:50];
  Mainzigotzufctzusync  MainzigotzufctzusyncR5 (gMainzigotzufctzusyncR5[18:0], callResR69);
  assign gMainzigotzunzucharzusyncR5 = gzdLLzicase63690[68:50];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR5 (gMainzigotzunzucharzusyncR5[18:0], callResR70);
  assign gMainzigotzutimezucodezusyncR5 = gzdLLzicase63690[68:50];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR5 (gMainzigotzutimezucodezusyncR5[18:0], callResR71);
  assign gReWireziPreludezizbzbR14 = {callResR70, callResR71};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR14 (gReWireziPreludezizbzbR14[1], gReWireziPreludezizbzbR14[0], callResR72);
  assign gReWireziPreludezizbzbR15 = {callResR69, callResR72};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR15 (gReWireziPreludezizbzbR15[1], gReWireziPreludezizbzbR15[0], callResR73);
  assign gzdLLzicase66593 = {callResR73, gzdLLzicase63690[49:25], gzdLLzicase63690[24:0]};
  assign gzdLLzicase63686 = {gzdLLzicase66593[49:25], gzdLLzicase66593[24:0]};
  assign gMainziautozustartzuzz1 = gzdLLzicase63686[49:25];
  Mainziautozustartzuzz1  Mainziautozustartzuzz1 (gMainziautozustartzuzz1[24:0], callResR74);
  assign gMainzigotzunullzusynczuregR2 = gzdLLzicase63686[49:25];
  Mainzigotzunullzusynczureg  MainzigotzunullzusynczuregR2 (gMainzigotzunullzusynczuregR2[24:0], callResR75);
  assign gReWireziPreludezizaza = {callResR74, callResR75};
  ReWireziPreludezizaza  ReWireziPreludezizaza (gReWireziPreludezizaza[1], gReWireziPreludezizaza[0], callResR76);
  assign gMainziautozustartzuzz1R1 = gzdLLzicase63686[49:25];
  Mainziautozustartzuzz1  Mainziautozustartzuzz1R1 (gMainziautozustartzuzz1R1[24:0], callResR77);
  assign gMainzigotzunullzusynczuregR3 = gzdLLzicase63686[49:25];
  Mainzigotzunullzusynczureg  MainzigotzunullzusynczuregR3 (gMainzigotzunullzusynczuregR3[24:0], callResR78);
  assign gReWireziPreludezizazaR1 = {callResR77, callResR78};
  ReWireziPreludezizaza  ReWireziPreludezizazaR1 (gReWireziPreludezizazaR1[1], gReWireziPreludezizazaR1[0], callResR79);
  assign gzdLLzicase66583 = {callResR79, gzdLLzicase63686[49:25], gzdLLzicase63686[24:0]};
  assign gzdLLzicase63683 = {gzdLLzicase66583[49:25], gzdLLzicase66583[24:0]};
  assign gMainzilinkzustartzuzz1 = gzdLLzicase63683[49:25];
  Mainzilinkzustartzuzz1  Mainzilinkzustartzuzz1 (gMainzilinkzustartzuzz1[24:0], callResR80);
  assign gMainzilinkzustartzuzz1R1 = gzdLLzicase63683[49:25];
  Mainzilinkzustartzuzz1  Mainzilinkzustartzuzz1R1 (gMainzilinkzustartzuzz1R1[24:0], callResR81);
  assign gzdLLzicase66573 = {callResR81, gzdLLzicase63683[24:0]};
  assign gzdLLzicase63680 = gzdLLzicase66573[24:0];
  assign gzdLLzilambda66566 = {gzdLLzicase63680[24:0], gzdLLzicase63680[24:0]};
  assign gzdLLzilambda63679 = gzdLLzilambda66566[49:0];
  assign gzdLLzicase63123R2 = gzdLLzilambda63679[49:25];
  zdLLzicase63123  zdLLzicase63123R2 (gzdLLzicase63123R2[24], gzdLLzicase63123R2[23], gzdLLzicase63123R2[22], gzdLLzicase63123R2[21], gzdLLzicase63123R2[20], gzdLLzicase63123R2[19], gzdLLzicase63123R2[18], gzdLLzicase63123R2[17], gzdLLzicase63123R2[16], gzdLLzicase63123R2[15], gzdLLzicase63123R2[14], gzdLLzicase63123R2[13], gzdLLzicase63123R2[12], gzdLLzicase63123R2[11], gzdLLzicase63123R2[10], gzdLLzicase63123R2[9], gzdLLzicase63123R2[8], gzdLLzicase63123R2[7], gzdLLzicase63123R2[6], gzdLLzicase63123R2[5], gzdLLzicase63123R2[4], gzdLLzicase63123R2[3], gzdLLzicase63123R2[2:0], callResR82);
  assign gzdLLzicase66575 = {callResR80, gzdLLzicase63683[24:0]};
  assign gzdLLzicase63681 = gzdLLzicase66575[24:0];
  assign gzdLLzilambda66571 = {gzdLLzicase63681[24:0], gzdLLzicase63681[24:0]};
  assign gzdLLzilambda63653 = gzdLLzilambda66571[49:0];
  assign gzdLLzicase63625 = gzdLLzilambda63653[49:25];
  zdLLzicase63625  zdLLzicase63625 (gzdLLzicase63625[24], gzdLLzicase63625[23], gzdLLzicase63625[22], gzdLLzicase63625[21], gzdLLzicase63625[20], gzdLLzicase63625[19], gzdLLzicase63625[18], gzdLLzicase63625[17], gzdLLzicase63625[16], gzdLLzicase63625[15], gzdLLzicase63625[14], gzdLLzicase63625[13], gzdLLzicase63625[12], gzdLLzicase63625[11], gzdLLzicase63625[10], gzdLLzicase63625[9], gzdLLzicase63625[8], gzdLLzicase63625[7], gzdLLzicase63625[6], gzdLLzicase63625[5], gzdLLzicase63625[4], gzdLLzicase63625[3], gzdLLzicase63625[2:0], callResR83);
  assign gzdLLzicase66585 = {callResR76, gzdLLzicase63686[24:0]};
  assign gzdLLzicase63684 = gzdLLzicase66585[24:0];
  assign gzdLLzilambda66580 = {gzdLLzicase63684[24:0], gzdLLzicase63684[24:0]};
  assign gzdLLzilambda63627 = gzdLLzilambda66580[49:0];
  assign gzdLLzicase63625R1 = gzdLLzilambda63627[49:25];
  zdLLzicase63625  zdLLzicase63625R1 (gzdLLzicase63625R1[24], gzdLLzicase63625R1[23], gzdLLzicase63625R1[22], gzdLLzicase63625R1[21], gzdLLzicase63625R1[20], gzdLLzicase63625R1[19], gzdLLzicase63625R1[18], gzdLLzicase63625R1[17], gzdLLzicase63625R1[16], gzdLLzicase63625R1[15], gzdLLzicase63625R1[14], gzdLLzicase63625R1[13], gzdLLzicase63625R1[12], gzdLLzicase63625R1[11], gzdLLzicase63625R1[10], gzdLLzicase63625R1[9], gzdLLzicase63625R1[8], gzdLLzicase63625R1[7], gzdLLzicase63625R1[6], gzdLLzicase63625R1[5], gzdLLzicase63625R1[4], gzdLLzicase63625R1[3], gzdLLzicase63625R1[2:0], callResR84);
  assign gzdLLzicase66595 = {callResR68, gzdLLzicase63690[24:0]};
  assign gzdLLzicase63687 = gzdLLzicase66595[24:0];
  assign gzdLLzilambda66590 = {gzdLLzicase63687[24:0], gzdLLzicase63687[24:0]};
  assign gzdLLzilambda63601 = gzdLLzilambda66590[49:0];
  assign gzdLLzicase63071R2 = gzdLLzilambda63601[49:25];
  zdLLzicase63071  zdLLzicase63071R2 (gzdLLzicase63071R2[24], gzdLLzicase63071R2[23], gzdLLzicase63071R2[22], gzdLLzicase63071R2[21], gzdLLzicase63071R2[20], gzdLLzicase63071R2[19], gzdLLzicase63071R2[18], gzdLLzicase63071R2[17], gzdLLzicase63071R2[16], gzdLLzicase63071R2[15], gzdLLzicase63071R2[14], gzdLLzicase63071R2[13], gzdLLzicase63071R2[12], gzdLLzicase63071R2[11], gzdLLzicase63071R2[10], gzdLLzicase63071R2[9], gzdLLzicase63071R2[8], gzdLLzicase63071R2[7], gzdLLzicase63071R2[6], gzdLLzicase63071R2[5], gzdLLzicase63071R2[4], gzdLLzicase63071R2[3], gzdLLzicase63071R2[2:0], callResR85);
  assign gzdLLzicase66985 = {callResR62, gzdLLzilambda63697[24:0]};
  assign gzdLLzicase63691 = gzdLLzicase66985[24:0];
  assign gzdLLzilambda66600 = {gzdLLzicase63691[24:0], gzdLLzicase63691[24:0]};
  assign gzdLLzilambda63575 = gzdLLzilambda66600[49:0];
  assign gzdLLzicase62993R6 = gzdLLzilambda63575[49:25];
  zdLLzicase62993  zdLLzicase62993R6 (gzdLLzicase62993R6[24], gzdLLzicase62993R6[23], gzdLLzicase62993R6[22], gzdLLzicase62993R6[21], gzdLLzicase62993R6[20], gzdLLzicase62993R6[19], gzdLLzicase62993R6[18], gzdLLzicase62993R6[17], gzdLLzicase62993R6[16], gzdLLzicase62993R6[15], gzdLLzicase62993R6[14], gzdLLzicase62993R6[13], gzdLLzicase62993R6[12], gzdLLzicase62993R6[11], gzdLLzicase62993R6[10], gzdLLzicase62993R6[9], gzdLLzicase62993R6[8], gzdLLzicase62993R6[7], gzdLLzicase62993R6[6], gzdLLzicase62993R6[5], gzdLLzicase62993R6[4], gzdLLzicase62993R6[3], gzdLLzicase62993R6[2:0], callResR86);
  assign gzdLLzilambda66979 = {gzdLLzilambda63697[68:50], (gzdLLzicase66985[25] == 1'h1) ? callResR86 : ((gzdLLzicase66595[25] == 1'h1) ? callResR85 : ((gzdLLzicase66585[25] == 1'h1) ? callResR84 : ((gzdLLzicase66575[25] == 1'h1) ? callResR83 : callResR82)))};
  assign gzdLLzicase66831R3 = {gzdLLzilambda66979[24:0], gzdLLzilambda66979[43:25]};
  zdLLzicase66831  zdLLzicase66831R3 (gzdLLzicase66831R3[43:19], gzdLLzicase66831R3[18:0], callResR87);
  assign gzdLLzilambda67458 = callResR87;
  assign gzdLLzicase67426R3 = gzdLLzilambda67458[39:0];
  zdLLzicase67426  zdLLzicase67426R3 (gzdLLzicase67426R3[39:25], gzdLLzicase67426R3[24:0], callResR88);
  assign gzdLLzilambda67453 = callResR88;
  assign gzdLLzicase67451 = gzdLLzilambda67453[44:0];
  assign gzdLLzilambda62531 = {gzdLLzicase67451[39:25], gzdLLzicase67451[24:0]};
  assign gzdLLzicase67553 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62553 = {gzdLLzicase67553[43:25], gzdLLzicase67553[24:0]};
  assign gMainzislsmzuerrorzuwait = {gzdLLzicase62553[43:25], gzdLLzicase62553[24:0]};
  assign gzdLLzilambda67377 = {gMainzislsmzuerrorzuwait[43:25], gMainzislsmzuerrorzuwait[24:0], gMainzislsmzuerrorzuwait[24:0]};
  assign gzdLLzicase67374 = {gzdLLzilambda67377[49:0], gzdLLzilambda67377[68:50]};
  assign gzdLLzilambda63497 = {gzdLLzicase67374[18:0], gzdLLzicase67374[68:44], gzdLLzicase67374[43:19]};
  assign gzdLLzicase63368 = gzdLLzilambda63497[49:25];
  assign gzdLLzilambda66972 = {gzdLLzilambda63497[68:50], {2'h2, gzdLLzicase63368[22], gzdLLzicase63368[21], 1'h0, gzdLLzicase63368[19], gzdLLzicase63368[18], gzdLLzicase63368[17], gzdLLzicase63368[16], gzdLLzicase63368[15], gzdLLzicase63368[14], gzdLLzicase63368[13], 1'h1, gzdLLzicase63368[11], gzdLLzicase63368[10], gzdLLzicase63368[9], gzdLLzicase63368[8], gzdLLzicase63368[7], gzdLLzicase63368[6], gzdLLzicase63368[5], gzdLLzicase63368[4], gzdLLzicase63368[3], gzdLLzicase63368[2:0]}};
  assign gzdLLzicase66969 = {gzdLLzilambda66972[24:0], gzdLLzilambda66972[43:25]};
  assign gzdLLzilambda63494 = {gzdLLzicase66969[18:0], gzdLLzicase66969[43:19]};
  assign gMainzigotzunullzusyncR4 = gzdLLzilambda63494[43:25];
  Mainzigotzunullzusync  MainzigotzunullzusyncR4 (gMainzigotzunullzusyncR4[18:0], callResR89);
  assign gMainzigotzunullzusyncR5 = gzdLLzilambda63494[43:25];
  Mainzigotzunullzusync  MainzigotzunullzusyncR5 (gMainzigotzunullzusyncR5[18:0], callResR90);
  assign idR2 = {callResR90, gzdLLzilambda63494[24:0]};
  assign gzdLLzicase66965 = {callResR89, gzdLLzilambda63494[24:0]};
  assign gzdLLzicase63396 = gzdLLzicase66965[24:0];
  assign gzdLLzilambda66532 = {gzdLLzicase63396[24:0], gzdLLzicase63396[24:0]};
  assign gzdLLzilambda63394 = gzdLLzilambda66532[49:0];
  assign gzdLLzicase63392R1 = gzdLLzilambda63394[49:25];
  zdLLzicase63392  zdLLzicase63392R1 (gzdLLzicase63392R1[24], gzdLLzicase63392R1[23], gzdLLzicase63392R1[22], gzdLLzicase63392R1[21], gzdLLzicase63392R1[20], gzdLLzicase63392R1[19], gzdLLzicase63392R1[18], gzdLLzicase63392R1[17], gzdLLzicase63392R1[16], gzdLLzicase63392R1[15], gzdLLzicase63392R1[14], gzdLLzicase63392R1[13], gzdLLzicase63392R1[12], gzdLLzicase63392R1[11], gzdLLzicase63392R1[10], gzdLLzicase63392R1[9], gzdLLzicase63392R1[8], gzdLLzicase63392R1[7], gzdLLzicase63392R1[6], gzdLLzicase63392R1[5], gzdLLzicase63392R1[4], gzdLLzicase63392R1[3], gzdLLzicase63392R1[2:0], callResR91);
  assign gzdLLzilambda66961 = {gzdLLzilambda63494[43:25], (gzdLLzicase66965[25] == 1'h1) ? callResR91 : idR2[24:0]};
  assign gzdLLzicase66958 = {gzdLLzilambda66961[24:0], gzdLLzilambda66961[43:25]};
  assign gzdLLzilambda63491 = {gzdLLzicase66958[18:0], gzdLLzicase66958[43:19]};
  assign gzdLLzilambda66954 = {gzdLLzilambda63491[43:25], gzdLLzilambda63491[24:0], gzdLLzilambda63491[24:0]};
  assign gzdLLzicase66951 = {gzdLLzilambda66954[49:0], gzdLLzilambda66954[68:50]};
  assign gzdLLzilambda63488 = {gzdLLzicase66951[18:0], gzdLLzicase66951[68:44], gzdLLzicase66951[43:19]};
  assign gMainzirxzuerrorzusyncR7 = gzdLLzilambda63488[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR7 (gMainzirxzuerrorzusyncR7[24:0], callResR92);
  assign gMainzirxzuerrorzusyncR8 = gzdLLzilambda63488[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR8 (gMainzirxzuerrorzusyncR8[24:0], callResR93);
  assign gzdLLzicase66945 = {callResR93, gzdLLzilambda63488[68:50], gzdLLzilambda63488[24:0]};
  assign gzdLLzicase63481 = {gzdLLzicase66945[43:25], gzdLLzicase66945[24:0]};
  assign gMainzigotzufctzusyncR6 = gzdLLzicase63481[43:25];
  Mainzigotzufctzusync  MainzigotzufctzusyncR6 (gMainzigotzufctzusyncR6[18:0], callResR94);
  assign gMainzigotzunzucharzusyncR6 = gzdLLzicase63481[43:25];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR6 (gMainzigotzunzucharzusyncR6[18:0], callResR95);
  assign gMainzigotzutimezucodezusyncR6 = gzdLLzicase63481[43:25];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR6 (gMainzigotzutimezucodezusyncR6[18:0], callResR96);
  assign gReWireziPreludezizbzbR16 = {callResR95, callResR96};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR16 (gReWireziPreludezizbzbR16[1], gReWireziPreludezizbzbR16[0], callResR97);
  assign gReWireziPreludezizbzbR17 = {callResR94, callResR97};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR17 (gReWireziPreludezizbzbR17[1], gReWireziPreludezizbzbR17[0], callResR98);
  assign gMainzigotzufctzusyncR7 = gzdLLzicase63481[43:25];
  Mainzigotzufctzusync  MainzigotzufctzusyncR7 (gMainzigotzufctzusyncR7[18:0], callResR99);
  assign gMainzigotzunzucharzusyncR7 = gzdLLzicase63481[43:25];
  Mainzigotzunzucharzusync  MainzigotzunzucharzusyncR7 (gMainzigotzunzucharzusyncR7[18:0], callResR100);
  assign gMainzigotzutimezucodezusyncR7 = gzdLLzicase63481[43:25];
  Mainzigotzutimezucodezusync  MainzigotzutimezucodezusyncR7 (gMainzigotzutimezucodezusyncR7[18:0], callResR101);
  assign gReWireziPreludezizbzbR18 = {callResR100, callResR101};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR18 (gReWireziPreludezizbzbR18[1], gReWireziPreludezizbzbR18[0], callResR102);
  assign gReWireziPreludezizbzbR19 = {callResR99, callResR102};
  ReWireziPreludezizbzb  ReWireziPreludezizbzbR19 (gReWireziPreludezizbzbR19[1], gReWireziPreludezizbzbR19[0], callResR103);
  assign gzdLLzicase66549 = {callResR103, gzdLLzicase63481[43:25], gzdLLzicase63481[24:0]};
  assign gzdLLzicase63478 = {gzdLLzicase66549[43:25], gzdLLzicase66549[24:0]};
  assign gMainziizuafterzu12p8zuusR4 = gzdLLzicase63478[43:25];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuusR4 (gMainziizuafterzu12p8zuusR4[18:0], callResR104);
  assign gMainziizuafterzu12p8zuusR5 = gzdLLzicase63478[43:25];
  Mainziizuafterzu12p8zuus  Mainziizuafterzu12p8zuusR5 (gMainziizuafterzu12p8zuusR5[18:0], callResR105);
  assign idR3 = {callResR105, gzdLLzicase63478[24:0]};
  assign gzdLLzicase66541 = {callResR104, gzdLLzicase63478[24:0]};
  assign gzdLLzicase63476 = gzdLLzicase66541[24:0];
  assign gzdLLzilambda66537 = {gzdLLzicase63476[24:0], gzdLLzicase63476[24:0]};
  assign gzdLLzilambda63474 = gzdLLzilambda66537[49:0];
  assign gzdLLzicase63472 = gzdLLzilambda63474[49:25];
  assign gzdLLzicase66551 = {callResR98, gzdLLzicase63481[24:0]};
  assign gzdLLzicase63479 = gzdLLzicase66551[24:0];
  assign gzdLLzilambda66546 = {gzdLLzicase63479[24:0], gzdLLzicase63479[24:0]};
  assign gzdLLzilambda63448 = gzdLLzilambda66546[49:0];
  assign gzdLLzicase63071R3 = gzdLLzilambda63448[49:25];
  zdLLzicase63071  zdLLzicase63071R3 (gzdLLzicase63071R3[24], gzdLLzicase63071R3[23], gzdLLzicase63071R3[22], gzdLLzicase63071R3[21], gzdLLzicase63071R3[20], gzdLLzicase63071R3[19], gzdLLzicase63071R3[18], gzdLLzicase63071R3[17], gzdLLzicase63071R3[16], gzdLLzicase63071R3[15], gzdLLzicase63071R3[14], gzdLLzicase63071R3[13], gzdLLzicase63071R3[12], gzdLLzicase63071R3[11], gzdLLzicase63071R3[10], gzdLLzicase63071R3[9], gzdLLzicase63071R3[8], gzdLLzicase63071R3[7], gzdLLzicase63071R3[6], gzdLLzicase63071R3[5], gzdLLzicase63071R3[4], gzdLLzicase63071R3[3], gzdLLzicase63071R3[2:0], callResR106);
  assign gzdLLzicase66947 = {callResR92, gzdLLzilambda63488[24:0]};
  assign gzdLLzicase63482 = gzdLLzicase66947[24:0];
  assign gzdLLzilambda66556 = {gzdLLzicase63482[24:0], gzdLLzicase63482[24:0]};
  assign gzdLLzilambda63422 = gzdLLzilambda66556[49:0];
  assign gzdLLzicase62993R7 = gzdLLzilambda63422[49:25];
  zdLLzicase62993  zdLLzicase62993R7 (gzdLLzicase62993R7[24], gzdLLzicase62993R7[23], gzdLLzicase62993R7[22], gzdLLzicase62993R7[21], gzdLLzicase62993R7[20], gzdLLzicase62993R7[19], gzdLLzicase62993R7[18], gzdLLzicase62993R7[17], gzdLLzicase62993R7[16], gzdLLzicase62993R7[15], gzdLLzicase62993R7[14], gzdLLzicase62993R7[13], gzdLLzicase62993R7[12], gzdLLzicase62993R7[11], gzdLLzicase62993R7[10], gzdLLzicase62993R7[9], gzdLLzicase62993R7[8], gzdLLzicase62993R7[7], gzdLLzicase62993R7[6], gzdLLzicase62993R7[5], gzdLLzicase62993R7[4], gzdLLzicase62993R7[3], gzdLLzicase62993R7[2:0], callResR107);
  assign gzdLLzilambda66942 = {gzdLLzilambda63488[68:50], (gzdLLzicase66947[25] == 1'h1) ? callResR107 : ((gzdLLzicase66551[25] == 1'h1) ? callResR106 : ((gzdLLzicase66541[25] == 1'h1) ? {gzdLLzicase63472[24], gzdLLzicase63472[23], gzdLLzicase63472[22], gzdLLzicase63472[21], gzdLLzicase63472[20], gzdLLzicase63472[19], gzdLLzicase63472[18], gzdLLzicase63472[17], gzdLLzicase63472[16], gzdLLzicase63472[15], gzdLLzicase63472[14], gzdLLzicase63472[13], gzdLLzicase63472[12], gzdLLzicase63472[11], gzdLLzicase63472[10], gzdLLzicase63472[9], gzdLLzicase63472[8], gzdLLzicase63472[7], gzdLLzicase63472[6], gzdLLzicase63472[5], gzdLLzicase63472[4], gzdLLzicase63472[3], 3'h2} : idR3[24:0]))};
  assign gzdLLzicase66831R4 = {gzdLLzilambda66942[24:0], gzdLLzilambda66942[43:25]};
  zdLLzicase66831  zdLLzicase66831R4 (gzdLLzicase66831R4[43:19], gzdLLzicase66831R4[18:0], callResR108);
  assign gzdLLzilambda67468 = callResR108;
  assign gzdLLzicase67426R4 = gzdLLzilambda67468[39:0];
  zdLLzicase67426  zdLLzicase67426R4 (gzdLLzicase67426R4[39:25], gzdLLzicase67426R4[24:0], callResR109);
  assign gzdLLzilambda67463 = callResR109;
  assign gzdLLzicase67461 = gzdLLzilambda67463[44:0];
  assign gzdLLzilambda62527 = {gzdLLzicase67461[39:25], gzdLLzicase67461[24:0]};
  assign gzdLLzicase67556 = {gzdLLzilambda62558[27:25], gzdLLzilambda62558[46:28], gzdLLzilambda62558[24:0]};
  assign gzdLLzicase62555 = {gzdLLzicase67556[43:25], gzdLLzicase67556[24:0]};
  assign gMainzislsmzuerrorzureset = {gzdLLzicase62555[43:25], gzdLLzicase62555[24:0]};
  assign gzdLLzilambda67365 = {gMainzislsmzuerrorzureset[43:25], gMainzislsmzuerrorzureset[24:0], gMainzislsmzuerrorzureset[24:0]};
  assign gzdLLzicase67362 = {gzdLLzilambda67365[49:0], gzdLLzilambda67365[68:50]};
  assign gzdLLzilambda63344 = {gzdLLzicase67362[18:0], gzdLLzicase67362[68:44], gzdLLzicase67362[43:19]};
  assign gzdLLzicase63176 = gzdLLzilambda63344[49:25];
  assign gzdLLzilambda66935 = {gzdLLzilambda63344[68:50], {gzdLLzicase63176[24], gzdLLzicase63176[23], 1'h0, gzdLLzicase63176[21], gzdLLzicase63176[20], gzdLLzicase63176[19], gzdLLzicase63176[18], gzdLLzicase63176[17], gzdLLzicase63176[16], 1'h0, gzdLLzicase63176[14], gzdLLzicase63176[13], gzdLLzicase63176[12], gzdLLzicase63176[11], gzdLLzicase63176[10], gzdLLzicase63176[9], gzdLLzicase63176[8], gzdLLzicase63176[7], gzdLLzicase63176[6], gzdLLzicase63176[5], gzdLLzicase63176[4], gzdLLzicase63176[3], gzdLLzicase63176[2:0]}};
  assign gzdLLzicase66932 = {gzdLLzilambda66935[24:0], gzdLLzilambda66935[43:25]};
  assign gzdLLzilambda63341 = {gzdLLzicase66932[18:0], gzdLLzicase66932[43:19]};
  assign gzdLLzilambda66928 = {gzdLLzilambda63341[43:25], gzdLLzilambda63341[24:0], gzdLLzilambda63341[24:0]};
  assign gzdLLzicase66925 = {gzdLLzilambda66928[49:0], gzdLLzilambda66928[68:50]};
  assign gzdLLzilambda63338 = {gzdLLzicase66925[18:0], gzdLLzicase66925[68:44], gzdLLzicase66925[43:19]};
  assign gzdLLzilambda66921 = {gzdLLzilambda63338[49:25], gzdLLzilambda63338[68:50], gzdLLzilambda63338[24:0], gzdLLzilambda63338[24:0]};
  assign gzdLLzicase66917 = {gzdLLzilambda66921[49:0], gzdLLzilambda66921[93:69], gzdLLzilambda66921[68:50]};
  assign gzdLLzilambda63335 = {gzdLLzicase66917[43:19], gzdLLzicase66917[18:0], gzdLLzicase66917[93:69], gzdLLzicase66917[68:44]};
  assign gzdLLzicase63201 = {gzdLLzilambda63335[49:25], gzdLLzilambda63335[93:69]};
  assign gMainzisendzutimezucodeR1 = gzdLLzicase63201[24:0];
  Mainzisendzutimezucode  MainzisendzutimezucodeR1 (gMainzisendzutimezucodeR1[24:0], callResR110);
  assign litR2 = callResR110;
  assign gzdLLzilambda66912 = {gzdLLzilambda63335[68:50], {gzdLLzicase63201[49], gzdLLzicase63201[48], gzdLLzicase63201[47], gzdLLzicase63201[46], gzdLLzicase63201[45], gzdLLzicase63201[44], gzdLLzicase63201[43], gzdLLzicase63201[42], gzdLLzicase63201[41], gzdLLzicase63201[40], (litR2[0] == 1'h1) ? 1'h1 : 1'h0, gzdLLzicase63201[38], gzdLLzicase63201[37], gzdLLzicase63201[36], gzdLLzicase63201[35], gzdLLzicase63201[34], gzdLLzicase63201[33], gzdLLzicase63201[32], gzdLLzicase63201[31], gzdLLzicase63201[30], gzdLLzicase63201[29], gzdLLzicase63201[28], gzdLLzicase63201[27:25]}};
  assign gzdLLzicase66909 = {gzdLLzilambda66912[24:0], gzdLLzilambda66912[43:25]};
  assign gzdLLzilambda63331 = {gzdLLzicase66909[18:0], gzdLLzicase66909[43:19]};
  assign gzdLLzilambda66905 = {gzdLLzilambda63331[43:25], gzdLLzilambda63331[24:0], gzdLLzilambda63331[24:0]};
  assign gzdLLzicase66902 = {gzdLLzilambda66905[49:0], gzdLLzilambda66905[68:50]};
  assign gzdLLzilambda63328 = {gzdLLzicase66902[18:0], gzdLLzicase66902[68:44], gzdLLzicase66902[43:19]};
  assign gMainzififozuavailablezuzz1 = gzdLLzilambda63328[49:25];
  Mainzififozuavailablezuzz1  Mainzififozuavailablezuzz1 (gMainzififozuavailablezuzz1[24:0], callResR111);
  assign gMainzififozuavailablezuzz1R1 = gzdLLzilambda63328[49:25];
  Mainzififozuavailablezuzz1  Mainzififozuavailablezuzz1R1 (gMainzififozuavailablezuzz1R1[24:0], callResR112);
  assign idR4 = {callResR112, gzdLLzilambda63328[24:0]};
  assign gzdLLzicase66898 = {callResR111, gzdLLzilambda63328[24:0]};
  assign gzdLLzicase63229 = gzdLLzicase66898[24:0];
  assign gzdLLzilambda66513 = {gzdLLzicase63229[24:0], gzdLLzicase63229[24:0]};
  assign gzdLLzilambda63227 = gzdLLzilambda66513[49:0];
  assign gzdLLzicase63225 = gzdLLzilambda63227[49:25];
  assign gzdLLzilambda66894 = {gzdLLzilambda63328[68:50], (gzdLLzicase66898[25] == 1'h1) ? {gzdLLzicase63225[24], gzdLLzicase63225[23], gzdLLzicase63225[22], 1'h0, gzdLLzicase63225[20], gzdLLzicase63225[19], gzdLLzicase63225[18], gzdLLzicase63225[17], gzdLLzicase63225[16], gzdLLzicase63225[15], gzdLLzicase63225[14], gzdLLzicase63225[13], gzdLLzicase63225[12], gzdLLzicase63225[11], gzdLLzicase63225[10], gzdLLzicase63225[9], gzdLLzicase63225[8], gzdLLzicase63225[7], gzdLLzicase63225[6], gzdLLzicase63225[5], gzdLLzicase63225[4], gzdLLzicase63225[3], gzdLLzicase63225[2:0]} : idR4[24:0]};
  assign gzdLLzicase66891 = {gzdLLzilambda66894[24:0], gzdLLzilambda66894[43:25]};
  assign gzdLLzilambda63325 = {gzdLLzicase66891[18:0], gzdLLzicase66891[43:19]};
  assign gzdLLzilambda66887 = {gzdLLzilambda63325[43:25], gzdLLzilambda63325[24:0], gzdLLzilambda63325[24:0]};
  assign gzdLLzicase66884 = {gzdLLzilambda66887[49:0], gzdLLzilambda66887[68:50]};
  assign gzdLLzilambda63322 = {gzdLLzicase66884[18:0], gzdLLzicase66884[68:44], gzdLLzicase66884[43:19]};
  assign gzdLLzicase63253 = gzdLLzilambda63322[49:25];
  assign gzdLLzilambda66880 = {gzdLLzilambda63322[68:50], {2'h0, gzdLLzicase63253[22], 1'h0, gzdLLzicase63253[20], 4'h0, gzdLLzicase63253[15], gzdLLzicase63253[14], gzdLLzicase63253[13], 1'h0, gzdLLzicase63253[11], gzdLLzicase63253[10], 1'h0, gzdLLzicase63253[8], gzdLLzicase63253[7], gzdLLzicase63253[6], gzdLLzicase63253[5], gzdLLzicase63253[4], gzdLLzicase63253[3], gzdLLzicase63253[2:0]}};
  assign gzdLLzicase66877 = {gzdLLzilambda66880[24:0], gzdLLzilambda66880[43:25]};
  assign gzdLLzilambda63319 = {gzdLLzicase66877[18:0], gzdLLzicase66877[43:19]};
  assign gzdLLzilambda66873 = {gzdLLzilambda63319[43:25], gzdLLzilambda63319[24:0], gzdLLzilambda63319[24:0]};
  assign gzdLLzicase66870 = {gzdLLzilambda66873[49:0], gzdLLzilambda66873[68:50]};
  assign gzdLLzilambda63316 = {gzdLLzicase66870[18:0], gzdLLzicase66870[68:44], gzdLLzicase66870[43:19]};
  assign gMainzirxzuerrorzusyncR9 = gzdLLzilambda63316[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR9 (gMainzirxzuerrorzusyncR9[24:0], callResR113);
  assign gMainzirxzuerrorzusyncR10 = gzdLLzilambda63316[49:25];
  Mainzirxzuerrorzusync  MainzirxzuerrorzusyncR10 (gMainzirxzuerrorzusyncR10[24:0], callResR114);
  assign gzdLLzicase66864 = {callResR114, gzdLLzilambda63316[68:50], gzdLLzilambda63316[24:0]};
  assign gzdLLzicase63309 = {gzdLLzicase66864[43:25], gzdLLzicase66864[24:0]};
  assign gMainziizuafterzu6p4zuus = gzdLLzicase63309[43:25];
  Mainziizuafterzu6p4zuus  Mainziizuafterzu6p4zuus (gMainziizuafterzu6p4zuus[18:0], callResR115);
  assign gMainziizuafterzu6p4zuusR1 = gzdLLzicase63309[43:25];
  Mainziizuafterzu6p4zuus  Mainziizuafterzu6p4zuusR1 (gMainziizuafterzu6p4zuusR1[18:0], callResR116);
  assign idR5 = {callResR116, gzdLLzicase63309[24:0]};
  assign gzdLLzicase66522 = {callResR115, gzdLLzicase63309[24:0]};
  assign gzdLLzicase63307 = gzdLLzicase66522[24:0];
  assign gzdLLzilambda66518 = {gzdLLzicase63307[24:0], gzdLLzicase63307[24:0]};
  assign gzdLLzilambda63305 = gzdLLzilambda66518[49:0];
  assign gzdLLzicase63303 = gzdLLzilambda63305[49:25];
  assign gzdLLzicase66866 = {callResR113, gzdLLzilambda63316[24:0]};
  assign gzdLLzicase63310 = gzdLLzicase66866[24:0];
  assign gzdLLzilambda66527 = {gzdLLzicase63310[24:0], gzdLLzicase63310[24:0]};
  assign gzdLLzilambda63279 = gzdLLzilambda66527[49:0];
  assign gzdLLzicase63123R3 = gzdLLzilambda63279[49:25];
  zdLLzicase63123  zdLLzicase63123R3 (gzdLLzicase63123R3[24], gzdLLzicase63123R3[23], gzdLLzicase63123R3[22], gzdLLzicase63123R3[21], gzdLLzicase63123R3[20], gzdLLzicase63123R3[19], gzdLLzicase63123R3[18], gzdLLzicase63123R3[17], gzdLLzicase63123R3[16], gzdLLzicase63123R3[15], gzdLLzicase63123R3[14], gzdLLzicase63123R3[13], gzdLLzicase63123R3[12], gzdLLzicase63123R3[11], gzdLLzicase63123R3[10], gzdLLzicase63123R3[9], gzdLLzicase63123R3[8], gzdLLzicase63123R3[7], gzdLLzicase63123R3[6], gzdLLzicase63123R3[5], gzdLLzicase63123R3[4], gzdLLzicase63123R3[3], gzdLLzicase63123R3[2:0], callResR117);
  assign gzdLLzilambda66861 = {gzdLLzilambda63316[68:50], (gzdLLzicase66866[25] == 1'h1) ? callResR117 : ((gzdLLzicase66522[25] == 1'h1) ? {gzdLLzicase63303[24], gzdLLzicase63303[23], gzdLLzicase63303[22], gzdLLzicase63303[21], 1'h1, gzdLLzicase63303[19], gzdLLzicase63303[18], gzdLLzicase63303[17], gzdLLzicase63303[16], gzdLLzicase63303[15], gzdLLzicase63303[14], gzdLLzicase63303[13], gzdLLzicase63303[12], gzdLLzicase63303[11], gzdLLzicase63303[10], gzdLLzicase63303[9], gzdLLzicase63303[8], gzdLLzicase63303[7], gzdLLzicase63303[6], gzdLLzicase63303[5], gzdLLzicase63303[4], gzdLLzicase63303[3], 3'h1} : idR5[24:0])};
  assign gzdLLzicase66831R5 = {gzdLLzilambda66861[24:0], gzdLLzilambda66861[43:25]};
  zdLLzicase66831  zdLLzicase66831R5 (gzdLLzicase66831R5[43:19], gzdLLzicase66831R5[18:0], callResR118);
  assign gzdLLzilambda67478 = callResR118;
  assign gzdLLzicase67426R5 = gzdLLzilambda67478[39:0];
  zdLLzicase67426  zdLLzicase67426R5 (gzdLLzicase67426R5[39:25], gzdLLzicase67426R5[24:0], callResR119);
  assign gzdLLzilambda67473 = callResR119;
  assign gzdLLzicase67471 = gzdLLzilambda67473[44:0];
  assign gzdLLzilambda62523 = {gzdLLzicase67471[39:25], gzdLLzicase67471[24:0]};
  assign res = (gzdLLzicase67556[46:44] == 3'h0) ? {1'h1, gzdLLzilambda62523[39:25], 4'h0, gzdLLzilambda62523[24:0]} : ((gzdLLzicase67553[46:44] == 3'h1) ? {1'h1, gzdLLzilambda62527[39:25], 4'h1, gzdLLzilambda62527[24:0]} : ((gzdLLzicase67550[46:44] == 3'h2) ? {1'h1, gzdLLzilambda62531[39:25], 4'h2, gzdLLzilambda62531[24:0]} : ((gzdLLzicase67547[46:44] == 3'h3) ? {1'h1, gzdLLzilambda62535[39:25], 4'h3, gzdLLzilambda62535[24:0]} : ((gzdLLzicase67544[46:44] == 3'h4) ? {1'h1, gzdLLzilambda62539[39:25], 4'h4, gzdLLzilambda62539[24:0]} : {1'h1, gzdLLzilambda62543[39:25], 4'h5, gzdLLzilambda62543[24:0]}))));
endmodule

module zdLLzicase66831 (input logic [24:0] arg0,
  input logic [18:0] arg1,
  output logic [39:0] res);
  logic [43:0] gMainzimkoutput;
  logic [68:0] gzdLLzilambda67341;
  logic [68:0] gzdLLzicase67338;
  logic [68:0] gzdLLzilambda62801;
  logic [24:0] gMainzitxzuen;
  logic [24:0] gzdLLzicase64167;
  logic [24:0] gMainzisendzunulls;
  logic [24:0] gzdLLzicase62921;
  logic [24:0] gMainzisendzufcts;
  logic [24:0] gzdLLzicase62873;
  logic [24:0] gMainzisendzunzuchar;
  logic [24:0] gzdLLzicase62897;
  logic [24:0] gMainzisendzutimezucode;
  logic [0:0] callRes;
  logic [24:0] gMainzirxzuen;
  logic [24:0] gzdLLzicase62825;
  logic [24:0] gMainzicharzusequencezuerror;
  logic [24:0] gzdLLzicase62517;
  logic [24:0] gMainzispacezuwirezuresetzunzuout;
  logic [24:0] gzdLLzicase64023;
  logic [24:0] gMainzitimerzu6p4zuuszureset;
  logic [24:0] gzdLLzicase64143;
  logic [24:0] gMainzitimerzu12p8zuuszustart;
  logic [24:0] gzdLLzicase64119;
  logic [24:0] gMainzistatzuinfozulinkzuupzutx;
  logic [24:0] gzdLLzicase64095;
  logic [24:0] gMainzistatzuinfozulinkzudownzutx;
  logic [24:0] gzdLLzicase64047;
  logic [24:0] gMainzistatzuinfozulinkzuupzuen;
  logic [24:0] gzdLLzicase64071;
  logic [18:0] gMainzigotzunullzusync;
  logic [0:0] callResR1;
  logic [18:0] gMainzigotzufctzusync;
  logic [0:0] callResR2;
  assign gMainzimkoutput = {arg1, arg0};
  assign gzdLLzilambda67341 = {gMainzimkoutput[43:25], gMainzimkoutput[24:0], gMainzimkoutput[24:0]};
  assign gzdLLzicase67338 = {gzdLLzilambda67341[49:0], gzdLLzilambda67341[68:50]};
  assign gzdLLzilambda62801 = {gzdLLzicase67338[18:0], gzdLLzicase67338[68:44], gzdLLzicase67338[43:19]};
  assign gMainzitxzuen = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64167 = gMainzitxzuen[24:0];
  assign gMainzisendzunulls = gzdLLzilambda62801[49:25];
  assign gzdLLzicase62921 = gMainzisendzunulls[24:0];
  assign gMainzisendzufcts = gzdLLzilambda62801[49:25];
  assign gzdLLzicase62873 = gMainzisendzufcts[24:0];
  assign gMainzisendzunzuchar = gzdLLzilambda62801[49:25];
  assign gzdLLzicase62897 = gMainzisendzunzuchar[24:0];
  assign gMainzisendzutimezucode = gzdLLzilambda62801[49:25];
  Mainzisendzutimezucode  Mainzisendzutimezucode (gMainzisendzutimezucode[24:0], callRes);
  assign gMainzirxzuen = gzdLLzilambda62801[49:25];
  assign gzdLLzicase62825 = gMainzirxzuen[24:0];
  assign gMainzicharzusequencezuerror = gzdLLzilambda62801[49:25];
  assign gzdLLzicase62517 = gMainzicharzusequencezuerror[24:0];
  assign gMainzispacezuwirezuresetzunzuout = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64023 = gMainzispacezuwirezuresetzunzuout[24:0];
  assign gMainzitimerzu6p4zuuszureset = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64143 = gMainzitimerzu6p4zuuszureset[24:0];
  assign gMainzitimerzu12p8zuuszustart = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64119 = gMainzitimerzu12p8zuuszustart[24:0];
  assign gMainzistatzuinfozulinkzuupzutx = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64095 = gMainzistatzuinfozulinkzuupzutx[24:0];
  assign gMainzistatzuinfozulinkzudownzutx = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64047 = gMainzistatzuinfozulinkzudownzutx[24:0];
  assign gMainzistatzuinfozulinkzuupzuen = gzdLLzilambda62801[49:25];
  assign gzdLLzicase64071 = gMainzistatzuinfozulinkzuupzuen[24:0];
  assign gMainzigotzunullzusync = gzdLLzilambda62801[68:50];
  Mainzigotzunullzusync  Mainzigotzunullzusync (gMainzigotzunullzusync[18:0], callResR1);
  assign gMainzigotzufctzusync = gzdLLzilambda62801[68:50];
  Mainzigotzufctzusync  Mainzigotzufctzusync (gMainzigotzufctzusync[18:0], callResR2);
  assign res = {gzdLLzicase64167[23], gzdLLzicase62921[18], gzdLLzicase62873[19], gzdLLzicase62897[17], callRes, gzdLLzicase62825[24], gzdLLzicase62517[9], gzdLLzicase64023[12], gzdLLzicase64143[21], gzdLLzicase64119[20], gzdLLzicase64095[13], gzdLLzicase64047[14], gzdLLzicase64071[15], callResR1, callResR2, gzdLLzilambda62801[24:0]};
endmodule

module zdLLzicase67426 (input logic [14:0] arg0,
  input logic [24:0] arg1,
  output logic [44:0] res);
  assign res = {5'h00, arg0, arg1};
endmodule

module Mainziautozustartzuzz1 (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62493;
  assign gzdLLzicase62493 = arg0;
  assign res = gzdLLzicase62493[7];
endmodule

module Mainzififozuavailablezuzz1 (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62582;
  assign gzdLLzicase62582 = arg0;
  assign res = gzdLLzicase62582[3];
endmodule

module Mainzigotzufctzusync (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62602;
  assign gzdLLzicase62602 = arg0;
  assign res = gzdLLzicase62602[2];
endmodule

module Mainzigotzunzucharzusync (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62622;
  assign gzdLLzicase62622 = arg0;
  assign res = gzdLLzicase62622[0];
endmodule

module Mainzigotzunullzusync (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62642;
  assign gzdLLzicase62642 = arg0;
  assign res = gzdLLzicase62642[3];
endmodule

module Mainzigotzunullzusynczureg (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62666;
  assign gzdLLzicase62666 = arg0;
  assign res = gzdLLzicase62666[22];
endmodule

module Mainzigotzutimezucodezusync (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62686;
  assign gzdLLzicase62686 = arg0;
  assign res = gzdLLzicase62686[1];
endmodule

module Mainziizuafterzu12p8zuus (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62706;
  assign gzdLLzicase62706 = arg0;
  assign res = gzdLLzicase62706[15];
endmodule

module Mainziizuafterzu6p4zuus (input logic [18:0] arg0,
  output logic [0:0] res);
  logic [18:0] gzdLLzicase62726;
  assign gzdLLzicase62726 = arg0;
  assign res = gzdLLzicase62726[14];
endmodule

module Mainzilinkzudisablezuzz1 (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62750;
  assign gzdLLzicase62750 = arg0;
  assign res = gzdLLzicase62750[11];
endmodule

module Mainzilinkzustartzuzz1 (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62774;
  assign gzdLLzicase62774 = arg0;
  assign res = gzdLLzicase62774[5];
endmodule

module Mainzirxzuerrorzusync (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62849;
  assign gzdLLzicase62849 = arg0;
  assign res = gzdLLzicase62849[10];
endmodule

module Mainzisendzutimezucode (input logic [24:0] arg0,
  output logic [0:0] res);
  logic [24:0] gzdLLzicase62945;
  assign gzdLLzicase62945 = arg0;
  assign res = gzdLLzicase62945[16];
endmodule

module ReWireziPreludezizaza (input logic [0:0] arg0,
  input logic [0:0] arg1,
  output logic [0:0] res);
  logic [1:0] lit;
  logic [1:0] id;
  assign lit = {arg0, arg1};
  assign id = {arg0, arg1};
  assign res = (id[1] == 1'h1) ? id[0] : 1'h0;
endmodule

module ReWireziPreludezizbzb (input logic [0:0] arg0,
  input logic [0:0] arg1,
  output logic [0:0] res);
  logic [1:0] id;
  logic [1:0] lit;
  assign id = {arg0, arg1};
  assign lit = {arg0, arg1};
  assign res = (lit[1] == 1'h1) ? 1'h1 : id[0];
endmodule